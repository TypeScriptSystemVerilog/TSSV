
  /* verilator lint_off DECLFILENAME */
  /* verilator lint_off UNUSED */
  
        

        
/* verilator lint_off WIDTH */        
module combN_tb 
   (
   input logic  clk,
   input logic  rst_b
   );

   logic [8:0] out;




endmodule
/* verilator lint_on WIDTH */        

