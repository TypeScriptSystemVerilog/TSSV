
        


interface AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION;

   logic [7:0] AWID;
   logic [47:0] AWADDR;
   logic [7:0] AWLEN;
   logic [2:0] AWSIZE;
   logic [1:0] AWBURST;
   logic  AWLOCK;
   logic [3:0] AWCACHE;
   logic [2:0] AWPROT;
   logic  AWVALID;
   logic  AWREADY;
   logic [127:0] WDATA;
   logic [15:0] WSTRB;
   logic  WLAST;
   logic  WVALID;
   logic  WREADY;
   logic [7:0] BID;
   logic [1:0] BRESP;
   logic  BVALID;
   logic  BREADY;
   logic [7:0] ARID;
   logic [47:0] ARADDR;
   logic [7:0] ARLEN;
   logic [2:0] ARSIZE;
   logic [1:0] ARBURST;
   logic  ARLOCK;
   logic [3:0] ARCACHE;
   logic [2:0] ARPROT;
   logic  ARVALID;
   logic  ARREADY;
   logic [7:0] RID;
   logic [127:0] RDATA;
   logic [1:0] RRESP;
   logic  RLAST;
   logic  RVALID;
   logic  RREADY;
   logic [3:0] ARQOS;
   logic [3:0] AWQOS;


    modport outward (
      output AWID,
      output AWADDR,
      output AWLEN,
      output AWSIZE,
      output AWBURST,
      output AWLOCK,
      output AWCACHE,
      output AWPROT,
      output AWQOS,
      output AWVALID,
      input AWREADY,
      output WDATA,
      output WSTRB,
      output WLAST,
      output WVALID,
      input WREADY,
      input BID,
      input BRESP,
      input BVALID,
      output BREADY,
      output ARID,
      output ARADDR,
      output ARLEN,
      output ARSIZE,
      output ARBURST,
      output ARLOCK,
      output ARCACHE,
      output ARPROT,
      output ARQOS,
      output ARVALID,
      input ARREADY,
      input RID,
      input RDATA,
      input RRESP,
      input RLAST,
      input RVALID,
      output RREADY
    );           

    modport inward (
      input AWID,
      input AWADDR,
      input AWLEN,
      input AWSIZE,
      input AWBURST,
      input AWLOCK,
      input AWCACHE,
      input AWPROT,
      input AWQOS,
      input AWVALID,
      output AWREADY,
      input WDATA,
      input WSTRB,
      input WLAST,
      input WVALID,
      output WREADY,
      output BID,
      output BRESP,
      output BVALID,
      input BREADY,
      input ARID,
      input ARADDR,
      input ARLEN,
      input ARSIZE,
      input ARBURST,
      input ARLOCK,
      input ARCACHE,
      input ARPROT,
      input ARQOS,
      input ARVALID,
      output ARREADY,
      output RID,
      output RDATA,
      output RRESP,
      output RLAST,
      output RVALID,
      input RREADY
    );           


endinterface
        
        
// Generated by CIRCT unknown git version

// Users can define 'STOP_COND' to add an extra gate to stop conditions.
`ifndef STOP_COND_
  `ifdef STOP_COND
    `define STOP_COND_ (`STOP_COND)
  `else  // STOP_COND
    `define STOP_COND_ 1
  `endif // STOP_COND
`endif // not def STOP_COND_

// Users can define 'ASSERT_VERBOSE_COND' to add an extra gate to assert error printing.
`ifndef ASSERT_VERBOSE_COND_
  `ifdef ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ (`ASSERT_VERBOSE_COND)
  `else  // ASSERT_VERBOSE_COND
    `define ASSERT_VERBOSE_COND_ 1
  `endif // ASSERT_VERBOSE_COND
`endif // not def ASSERT_VERBOSE_COND_

// Include register initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS


// Include rmemory initializers in init blocks unless synthesis is set
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

// Standard header to adapt well known macros for register randomization.

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_
module AXI4XBar2x4_inner(
  input          clock,
                 reset,
  output         master1_aw_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master1_aw_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master1_aw_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [47:0]  master1_aw_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master1_aw_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master1_aw_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [1:0]   master1_aw_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master1_aw_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master1_aw_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master1_aw_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master1_aw_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master1_w_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master1_w_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [127:0] master1_w_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [15:0]  master1_w_bits_strb,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master1_w_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:64:9
                 master1_b_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master1_b_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [7:0]   master1_b_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [1:0]   master1_b_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master1_ar_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master1_ar_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master1_ar_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [47:0]  master1_ar_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master1_ar_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master1_ar_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [1:0]   master1_ar_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master1_ar_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master1_ar_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master1_ar_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master1_ar_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master1_r_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master1_r_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [7:0]   master1_r_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [127:0] master1_r_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [1:0]   master1_r_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master1_r_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:64:9
                 master2_aw_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master2_aw_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master2_aw_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [47:0]  master2_aw_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master2_aw_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master2_aw_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [1:0]   master2_aw_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master2_aw_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master2_aw_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master2_aw_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master2_aw_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master2_w_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master2_w_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [127:0] master2_w_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [15:0]  master2_w_bits_strb,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master2_w_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:64:9
                 master2_b_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master2_b_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [7:0]   master2_b_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [1:0]   master2_b_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master2_ar_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master2_ar_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master2_ar_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [47:0]  master2_ar_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [7:0]   master2_ar_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master2_ar_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [1:0]   master2_ar_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master2_ar_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master2_ar_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [2:0]   master2_ar_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input  [3:0]   master2_ar_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          master2_r_ready,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master2_r_valid,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [7:0]   master2_r_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [127:0] master2_r_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output [1:0]   master2_r_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  output         master2_r_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:64:9
  input          slave1_aw_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave1_aw_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave1_aw_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave1_aw_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave1_aw_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave1_aw_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave1_aw_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave1_aw_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave1_aw_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave1_aw_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave1_aw_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave1_w_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave1_w_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [127:0] slave1_w_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [15:0]  slave1_w_bits_strb,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave1_w_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:67:9
                 slave1_b_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave1_b_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave1_b_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave1_b_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave1_ar_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave1_ar_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave1_ar_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave1_ar_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave1_ar_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave1_ar_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave1_ar_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave1_ar_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave1_ar_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave1_ar_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave1_ar_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave1_r_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave1_r_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave1_r_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [127:0] slave1_r_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave1_r_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave1_r_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:67:9
                 slave2_aw_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave2_aw_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave2_aw_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave2_aw_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave2_aw_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave2_aw_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave2_aw_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave2_aw_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave2_aw_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave2_aw_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave2_aw_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave2_w_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave2_w_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [127:0] slave2_w_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [15:0]  slave2_w_bits_strb,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave2_w_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:67:9
                 slave2_b_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave2_b_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave2_b_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave2_b_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave2_ar_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave2_ar_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave2_ar_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave2_ar_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave2_ar_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave2_ar_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave2_ar_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave2_ar_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave2_ar_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave2_ar_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave2_ar_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave2_r_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave2_r_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave2_r_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [127:0] slave2_r_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave2_r_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave2_r_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:67:9
                 slave3_aw_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave3_aw_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave3_aw_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave3_aw_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave3_aw_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave3_aw_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave3_aw_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave3_aw_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave3_aw_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave3_aw_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave3_aw_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave3_w_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave3_w_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [127:0] slave3_w_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [15:0]  slave3_w_bits_strb,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave3_w_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:67:9
                 slave3_b_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave3_b_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave3_b_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave3_b_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave3_ar_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave3_ar_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave3_ar_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave3_ar_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave3_ar_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave3_ar_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave3_ar_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave3_ar_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave3_ar_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave3_ar_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave3_ar_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave3_r_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave3_r_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave3_r_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [127:0] slave3_r_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave3_r_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave3_r_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:67:9
                 slave4_aw_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave4_aw_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave4_aw_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave4_aw_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave4_aw_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave4_aw_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave4_aw_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave4_aw_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave4_aw_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave4_aw_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave4_aw_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave4_w_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave4_w_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [127:0] slave4_w_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [15:0]  slave4_w_bits_strb,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave4_w_bits_last,	// src/main/scala/componentgen/componentgenModule.scala:67:9
                 slave4_b_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave4_b_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave4_b_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave4_b_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave4_ar_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave4_ar_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave4_ar_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [47:0]  slave4_ar_bits_addr,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [7:0]   slave4_ar_bits_len,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave4_ar_bits_size,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [1:0]   slave4_ar_bits_burst,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave4_ar_bits_lock,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave4_ar_bits_cache,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [2:0]   slave4_ar_bits_prot,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output [3:0]   slave4_ar_bits_qos,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  output         slave4_r_ready,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave4_r_valid,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [7:0]   slave4_r_bits_id,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [127:0] slave4_r_bits_data,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input  [1:0]   slave4_r_bits_resp,	// src/main/scala/componentgen/componentgenModule.scala:67:9
  input          slave4_r_bits_last	// src/main/scala/componentgen/componentgenModule.scala:67:9
);

  wire [2:0]   xbar_in_1_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_1_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_0_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_0_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_auto_anon_out_3_r_bits_last;
  wire [1:0]   xbar_auto_anon_out_3_r_bits_resp;
  wire [127:0] xbar_auto_anon_out_3_r_bits_data;
  wire [2:0]   xbar_auto_anon_out_3_r_bits_id;
  wire         xbar_auto_anon_out_3_r_valid;
  wire         xbar_auto_anon_out_3_r_ready;
  wire [3:0]   xbar_auto_anon_out_3_ar_bits_qos;
  wire [2:0]   xbar_auto_anon_out_3_ar_bits_prot;
  wire [3:0]   xbar_auto_anon_out_3_ar_bits_cache;
  wire         xbar_auto_anon_out_3_ar_bits_lock;
  wire [1:0]   xbar_auto_anon_out_3_ar_bits_burst;
  wire [2:0]   xbar_auto_anon_out_3_ar_bits_size;
  wire [7:0]   xbar_auto_anon_out_3_ar_bits_len;
  wire [29:0]  xbar_auto_anon_out_3_ar_bits_addr;
  wire [2:0]   xbar_auto_anon_out_3_ar_bits_id;
  wire         xbar_auto_anon_out_3_ar_valid;
  wire         xbar_auto_anon_out_3_ar_ready;
  wire [1:0]   xbar_auto_anon_out_3_b_bits_resp;
  wire [2:0]   xbar_auto_anon_out_3_b_bits_id;
  wire         xbar_auto_anon_out_3_b_valid;
  wire         xbar_auto_anon_out_3_b_ready;
  wire         xbar_auto_anon_out_3_w_bits_last;
  wire [15:0]  xbar_auto_anon_out_3_w_bits_strb;
  wire [127:0] xbar_auto_anon_out_3_w_bits_data;
  wire         xbar_auto_anon_out_3_w_valid;
  wire         xbar_auto_anon_out_3_w_ready;
  wire [3:0]   xbar_auto_anon_out_3_aw_bits_qos;
  wire [2:0]   xbar_auto_anon_out_3_aw_bits_prot;
  wire [3:0]   xbar_auto_anon_out_3_aw_bits_cache;
  wire         xbar_auto_anon_out_3_aw_bits_lock;
  wire [1:0]   xbar_auto_anon_out_3_aw_bits_burst;
  wire [2:0]   xbar_auto_anon_out_3_aw_bits_size;
  wire [7:0]   xbar_auto_anon_out_3_aw_bits_len;
  wire [29:0]  xbar_auto_anon_out_3_aw_bits_addr;
  wire [2:0]   xbar_auto_anon_out_3_aw_bits_id;
  wire         xbar_auto_anon_out_3_aw_valid;
  wire         xbar_auto_anon_out_3_aw_ready;
  wire         xbar_auto_anon_out_2_r_bits_last;
  wire [1:0]   xbar_auto_anon_out_2_r_bits_resp;
  wire [127:0] xbar_auto_anon_out_2_r_bits_data;
  wire [2:0]   xbar_auto_anon_out_2_r_bits_id;
  wire         xbar_auto_anon_out_2_r_valid;
  wire         xbar_auto_anon_out_2_r_ready;
  wire [3:0]   xbar_auto_anon_out_2_ar_bits_qos;
  wire [2:0]   xbar_auto_anon_out_2_ar_bits_prot;
  wire [3:0]   xbar_auto_anon_out_2_ar_bits_cache;
  wire         xbar_auto_anon_out_2_ar_bits_lock;
  wire [1:0]   xbar_auto_anon_out_2_ar_bits_burst;
  wire [2:0]   xbar_auto_anon_out_2_ar_bits_size;
  wire [7:0]   xbar_auto_anon_out_2_ar_bits_len;
  wire [29:0]  xbar_auto_anon_out_2_ar_bits_addr;
  wire [2:0]   xbar_auto_anon_out_2_ar_bits_id;
  wire         xbar_auto_anon_out_2_ar_valid;
  wire         xbar_auto_anon_out_2_ar_ready;
  wire [1:0]   xbar_auto_anon_out_2_b_bits_resp;
  wire [2:0]   xbar_auto_anon_out_2_b_bits_id;
  wire         xbar_auto_anon_out_2_b_valid;
  wire         xbar_auto_anon_out_2_b_ready;
  wire         xbar_auto_anon_out_2_w_bits_last;
  wire [15:0]  xbar_auto_anon_out_2_w_bits_strb;
  wire [127:0] xbar_auto_anon_out_2_w_bits_data;
  wire         xbar_auto_anon_out_2_w_valid;
  wire         xbar_auto_anon_out_2_w_ready;
  wire [3:0]   xbar_auto_anon_out_2_aw_bits_qos;
  wire [2:0]   xbar_auto_anon_out_2_aw_bits_prot;
  wire [3:0]   xbar_auto_anon_out_2_aw_bits_cache;
  wire         xbar_auto_anon_out_2_aw_bits_lock;
  wire [1:0]   xbar_auto_anon_out_2_aw_bits_burst;
  wire [2:0]   xbar_auto_anon_out_2_aw_bits_size;
  wire [7:0]   xbar_auto_anon_out_2_aw_bits_len;
  wire [29:0]  xbar_auto_anon_out_2_aw_bits_addr;
  wire [2:0]   xbar_auto_anon_out_2_aw_bits_id;
  wire         xbar_auto_anon_out_2_aw_valid;
  wire         xbar_auto_anon_out_2_aw_ready;
  wire         xbar_auto_anon_out_1_r_bits_last;
  wire [1:0]   xbar_auto_anon_out_1_r_bits_resp;
  wire [127:0] xbar_auto_anon_out_1_r_bits_data;
  wire [2:0]   xbar_auto_anon_out_1_r_bits_id;
  wire         xbar_auto_anon_out_1_r_valid;
  wire         xbar_auto_anon_out_1_r_ready;
  wire [3:0]   xbar_auto_anon_out_1_ar_bits_qos;
  wire [2:0]   xbar_auto_anon_out_1_ar_bits_prot;
  wire [3:0]   xbar_auto_anon_out_1_ar_bits_cache;
  wire         xbar_auto_anon_out_1_ar_bits_lock;
  wire [1:0]   xbar_auto_anon_out_1_ar_bits_burst;
  wire [2:0]   xbar_auto_anon_out_1_ar_bits_size;
  wire [7:0]   xbar_auto_anon_out_1_ar_bits_len;
  wire [28:0]  xbar_auto_anon_out_1_ar_bits_addr;
  wire [2:0]   xbar_auto_anon_out_1_ar_bits_id;
  wire         xbar_auto_anon_out_1_ar_valid;
  wire         xbar_auto_anon_out_1_ar_ready;
  wire [1:0]   xbar_auto_anon_out_1_b_bits_resp;
  wire [2:0]   xbar_auto_anon_out_1_b_bits_id;
  wire         xbar_auto_anon_out_1_b_valid;
  wire         xbar_auto_anon_out_1_b_ready;
  wire         xbar_auto_anon_out_1_w_bits_last;
  wire [15:0]  xbar_auto_anon_out_1_w_bits_strb;
  wire [127:0] xbar_auto_anon_out_1_w_bits_data;
  wire         xbar_auto_anon_out_1_w_valid;
  wire         xbar_auto_anon_out_1_w_ready;
  wire [3:0]   xbar_auto_anon_out_1_aw_bits_qos;
  wire [2:0]   xbar_auto_anon_out_1_aw_bits_prot;
  wire [3:0]   xbar_auto_anon_out_1_aw_bits_cache;
  wire         xbar_auto_anon_out_1_aw_bits_lock;
  wire [1:0]   xbar_auto_anon_out_1_aw_bits_burst;
  wire [2:0]   xbar_auto_anon_out_1_aw_bits_size;
  wire [7:0]   xbar_auto_anon_out_1_aw_bits_len;
  wire [28:0]  xbar_auto_anon_out_1_aw_bits_addr;
  wire [2:0]   xbar_auto_anon_out_1_aw_bits_id;
  wire         xbar_auto_anon_out_1_aw_valid;
  wire         xbar_auto_anon_out_1_aw_ready;
  wire         xbar_auto_anon_out_0_r_bits_last;
  wire [1:0]   xbar_auto_anon_out_0_r_bits_resp;
  wire [127:0] xbar_auto_anon_out_0_r_bits_data;
  wire [2:0]   xbar_auto_anon_out_0_r_bits_id;
  wire         xbar_auto_anon_out_0_r_valid;
  wire         xbar_auto_anon_out_0_r_ready;
  wire [3:0]   xbar_auto_anon_out_0_ar_bits_qos;
  wire [2:0]   xbar_auto_anon_out_0_ar_bits_prot;
  wire [3:0]   xbar_auto_anon_out_0_ar_bits_cache;
  wire         xbar_auto_anon_out_0_ar_bits_lock;
  wire [1:0]   xbar_auto_anon_out_0_ar_bits_burst;
  wire [2:0]   xbar_auto_anon_out_0_ar_bits_size;
  wire [7:0]   xbar_auto_anon_out_0_ar_bits_len;
  wire [27:0]  xbar_auto_anon_out_0_ar_bits_addr;
  wire [2:0]   xbar_auto_anon_out_0_ar_bits_id;
  wire         xbar_auto_anon_out_0_ar_valid;
  wire         xbar_auto_anon_out_0_ar_ready;
  wire [1:0]   xbar_auto_anon_out_0_b_bits_resp;
  wire [2:0]   xbar_auto_anon_out_0_b_bits_id;
  wire         xbar_auto_anon_out_0_b_valid;
  wire         xbar_auto_anon_out_0_b_ready;
  wire         xbar_auto_anon_out_0_w_bits_last;
  wire [15:0]  xbar_auto_anon_out_0_w_bits_strb;
  wire [127:0] xbar_auto_anon_out_0_w_bits_data;
  wire         xbar_auto_anon_out_0_w_valid;
  wire         xbar_auto_anon_out_0_w_ready;
  wire [3:0]   xbar_auto_anon_out_0_aw_bits_qos;
  wire [2:0]   xbar_auto_anon_out_0_aw_bits_prot;
  wire [3:0]   xbar_auto_anon_out_0_aw_bits_cache;
  wire         xbar_auto_anon_out_0_aw_bits_lock;
  wire [1:0]   xbar_auto_anon_out_0_aw_bits_burst;
  wire [2:0]   xbar_auto_anon_out_0_aw_bits_size;
  wire [7:0]   xbar_auto_anon_out_0_aw_bits_len;
  wire [27:0]  xbar_auto_anon_out_0_aw_bits_addr;
  wire [2:0]   xbar_auto_anon_out_0_aw_bits_id;
  wire         xbar_auto_anon_out_0_aw_valid;
  wire         xbar_auto_anon_out_0_aw_ready;
  wire         xbar_auto_anon_in_1_r_bits_last;
  wire [1:0]   xbar_auto_anon_in_1_r_bits_resp;
  wire [127:0] xbar_auto_anon_in_1_r_bits_data;
  wire [1:0]   xbar_auto_anon_in_1_r_bits_id;
  wire         xbar_auto_anon_in_1_r_valid;
  wire         xbar_auto_anon_in_1_r_ready;
  wire [3:0]   xbar_auto_anon_in_1_ar_bits_qos;
  wire [2:0]   xbar_auto_anon_in_1_ar_bits_prot;
  wire [3:0]   xbar_auto_anon_in_1_ar_bits_cache;
  wire         xbar_auto_anon_in_1_ar_bits_lock;
  wire [1:0]   xbar_auto_anon_in_1_ar_bits_burst;
  wire [2:0]   xbar_auto_anon_in_1_ar_bits_size;
  wire [7:0]   xbar_auto_anon_in_1_ar_bits_len;
  wire [29:0]  xbar_auto_anon_in_1_ar_bits_addr;
  wire [1:0]   xbar_auto_anon_in_1_ar_bits_id;
  wire         xbar_auto_anon_in_1_ar_valid;
  wire         xbar_auto_anon_in_1_ar_ready;
  wire [1:0]   xbar_auto_anon_in_1_b_bits_resp;
  wire [1:0]   xbar_auto_anon_in_1_b_bits_id;
  wire         xbar_auto_anon_in_1_b_valid;
  wire         xbar_auto_anon_in_1_b_ready;
  wire         xbar_auto_anon_in_1_w_bits_last;
  wire [15:0]  xbar_auto_anon_in_1_w_bits_strb;
  wire [127:0] xbar_auto_anon_in_1_w_bits_data;
  wire         xbar_auto_anon_in_1_w_valid;
  wire         xbar_auto_anon_in_1_w_ready;
  wire [3:0]   xbar_auto_anon_in_1_aw_bits_qos;
  wire [2:0]   xbar_auto_anon_in_1_aw_bits_prot;
  wire [3:0]   xbar_auto_anon_in_1_aw_bits_cache;
  wire         xbar_auto_anon_in_1_aw_bits_lock;
  wire [1:0]   xbar_auto_anon_in_1_aw_bits_burst;
  wire [2:0]   xbar_auto_anon_in_1_aw_bits_size;
  wire [7:0]   xbar_auto_anon_in_1_aw_bits_len;
  wire [29:0]  xbar_auto_anon_in_1_aw_bits_addr;
  wire [1:0]   xbar_auto_anon_in_1_aw_bits_id;
  wire         xbar_auto_anon_in_1_aw_valid;
  wire         xbar_auto_anon_in_1_aw_ready;
  wire         xbar_auto_anon_in_0_r_bits_last;
  wire [1:0]   xbar_auto_anon_in_0_r_bits_resp;
  wire [127:0] xbar_auto_anon_in_0_r_bits_data;
  wire         xbar_auto_anon_in_0_r_valid;
  wire         xbar_auto_anon_in_0_r_ready;
  wire [3:0]   xbar_auto_anon_in_0_ar_bits_qos;
  wire [2:0]   xbar_auto_anon_in_0_ar_bits_prot;
  wire [3:0]   xbar_auto_anon_in_0_ar_bits_cache;
  wire         xbar_auto_anon_in_0_ar_bits_lock;
  wire [1:0]   xbar_auto_anon_in_0_ar_bits_burst;
  wire [2:0]   xbar_auto_anon_in_0_ar_bits_size;
  wire [7:0]   xbar_auto_anon_in_0_ar_bits_len;
  wire [29:0]  xbar_auto_anon_in_0_ar_bits_addr;
  wire         xbar_auto_anon_in_0_ar_bits_id;
  wire         xbar_auto_anon_in_0_ar_valid;
  wire         xbar_auto_anon_in_0_ar_ready;
  wire [1:0]   xbar_auto_anon_in_0_b_bits_resp;
  wire         xbar_auto_anon_in_0_b_valid;
  wire         xbar_auto_anon_in_0_b_ready;
  wire         xbar_auto_anon_in_0_w_bits_last;
  wire [15:0]  xbar_auto_anon_in_0_w_bits_strb;
  wire [127:0] xbar_auto_anon_in_0_w_bits_data;
  wire         xbar_auto_anon_in_0_w_valid;
  wire         xbar_auto_anon_in_0_w_ready;
  wire [3:0]   xbar_auto_anon_in_0_aw_bits_qos;
  wire [2:0]   xbar_auto_anon_in_0_aw_bits_prot;
  wire [3:0]   xbar_auto_anon_in_0_aw_bits_cache;
  wire         xbar_auto_anon_in_0_aw_bits_lock;
  wire [1:0]   xbar_auto_anon_in_0_aw_bits_burst;
  wire [2:0]   xbar_auto_anon_in_0_aw_bits_size;
  wire [7:0]   xbar_auto_anon_in_0_aw_bits_len;
  wire [29:0]  xbar_auto_anon_in_0_aw_bits_addr;
  wire         xbar_auto_anon_in_0_aw_bits_id;
  wire         xbar_auto_anon_in_0_aw_valid;
  wire         xbar_auto_anon_in_0_aw_ready;
  wire [1:0]   _ram_ext_R0_data;	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  wire [1:0]   _ram_ext_R0_data_0;	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  wire [1:0]   _ram_ext_R0_data_1;	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  wire [1:0]   _ram_ext_R0_data_2;	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  wire [3:0]   _ram_ext_R0_data_3;	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  wire [3:0]   _ram_ext_R0_data_4;	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  wire         master1_aw_valid_0 = master1_aw_valid;
  wire [7:0]   master1_aw_bits_id_0 = master1_aw_bits_id;
  wire [47:0]  master1_aw_bits_addr_0 = master1_aw_bits_addr;
  wire [7:0]   master1_aw_bits_len_0 = master1_aw_bits_len;
  wire [2:0]   master1_aw_bits_size_0 = master1_aw_bits_size;
  wire [1:0]   master1_aw_bits_burst_0 = master1_aw_bits_burst;
  wire         master1_aw_bits_lock_0 = master1_aw_bits_lock;
  wire [3:0]   master1_aw_bits_cache_0 = master1_aw_bits_cache;
  wire [2:0]   master1_aw_bits_prot_0 = master1_aw_bits_prot;
  wire [3:0]   master1_aw_bits_qos_0 = master1_aw_bits_qos;
  wire         master1_w_valid_0 = master1_w_valid;
  wire [127:0] master1_w_bits_data_0 = master1_w_bits_data;
  wire [15:0]  master1_w_bits_strb_0 = master1_w_bits_strb;
  wire         master1_w_bits_last_0 = master1_w_bits_last;
  wire         master1_b_ready_0 = master1_b_ready;
  wire         master1_ar_valid_0 = master1_ar_valid;
  wire [7:0]   master1_ar_bits_id_0 = master1_ar_bits_id;
  wire [47:0]  master1_ar_bits_addr_0 = master1_ar_bits_addr;
  wire [7:0]   master1_ar_bits_len_0 = master1_ar_bits_len;
  wire [2:0]   master1_ar_bits_size_0 = master1_ar_bits_size;
  wire [1:0]   master1_ar_bits_burst_0 = master1_ar_bits_burst;
  wire         master1_ar_bits_lock_0 = master1_ar_bits_lock;
  wire [3:0]   master1_ar_bits_cache_0 = master1_ar_bits_cache;
  wire [2:0]   master1_ar_bits_prot_0 = master1_ar_bits_prot;
  wire [3:0]   master1_ar_bits_qos_0 = master1_ar_bits_qos;
  wire         master1_r_ready_0 = master1_r_ready;
  wire         master2_aw_valid_0 = master2_aw_valid;
  wire [7:0]   master2_aw_bits_id_0 = master2_aw_bits_id;
  wire [47:0]  master2_aw_bits_addr_0 = master2_aw_bits_addr;
  wire [7:0]   master2_aw_bits_len_0 = master2_aw_bits_len;
  wire [2:0]   master2_aw_bits_size_0 = master2_aw_bits_size;
  wire [1:0]   master2_aw_bits_burst_0 = master2_aw_bits_burst;
  wire         master2_aw_bits_lock_0 = master2_aw_bits_lock;
  wire [3:0]   master2_aw_bits_cache_0 = master2_aw_bits_cache;
  wire [2:0]   master2_aw_bits_prot_0 = master2_aw_bits_prot;
  wire [3:0]   master2_aw_bits_qos_0 = master2_aw_bits_qos;
  wire         master2_w_valid_0 = master2_w_valid;
  wire [127:0] master2_w_bits_data_0 = master2_w_bits_data;
  wire [15:0]  master2_w_bits_strb_0 = master2_w_bits_strb;
  wire         master2_w_bits_last_0 = master2_w_bits_last;
  wire         master2_b_ready_0 = master2_b_ready;
  wire         master2_ar_valid_0 = master2_ar_valid;
  wire [7:0]   master2_ar_bits_id_0 = master2_ar_bits_id;
  wire [47:0]  master2_ar_bits_addr_0 = master2_ar_bits_addr;
  wire [7:0]   master2_ar_bits_len_0 = master2_ar_bits_len;
  wire [2:0]   master2_ar_bits_size_0 = master2_ar_bits_size;
  wire [1:0]   master2_ar_bits_burst_0 = master2_ar_bits_burst;
  wire         master2_ar_bits_lock_0 = master2_ar_bits_lock;
  wire [3:0]   master2_ar_bits_cache_0 = master2_ar_bits_cache;
  wire [2:0]   master2_ar_bits_prot_0 = master2_ar_bits_prot;
  wire [3:0]   master2_ar_bits_qos_0 = master2_ar_bits_qos;
  wire         master2_r_ready_0 = master2_r_ready;
  wire         slave1_aw_ready_0 = slave1_aw_ready;
  wire         slave1_w_ready_0 = slave1_w_ready;
  wire         slave1_b_valid_0 = slave1_b_valid;
  wire [7:0]   slave1_b_bits_id_0 = slave1_b_bits_id;
  wire [1:0]   slave1_b_bits_resp_0 = slave1_b_bits_resp;
  wire         slave1_ar_ready_0 = slave1_ar_ready;
  wire         slave1_r_valid_0 = slave1_r_valid;
  wire [7:0]   slave1_r_bits_id_0 = slave1_r_bits_id;
  wire [127:0] slave1_r_bits_data_0 = slave1_r_bits_data;
  wire [1:0]   slave1_r_bits_resp_0 = slave1_r_bits_resp;
  wire         slave1_r_bits_last_0 = slave1_r_bits_last;
  wire         slave2_aw_ready_0 = slave2_aw_ready;
  wire         slave2_w_ready_0 = slave2_w_ready;
  wire         slave2_b_valid_0 = slave2_b_valid;
  wire [7:0]   slave2_b_bits_id_0 = slave2_b_bits_id;
  wire [1:0]   slave2_b_bits_resp_0 = slave2_b_bits_resp;
  wire         slave2_ar_ready_0 = slave2_ar_ready;
  wire         slave2_r_valid_0 = slave2_r_valid;
  wire [7:0]   slave2_r_bits_id_0 = slave2_r_bits_id;
  wire [127:0] slave2_r_bits_data_0 = slave2_r_bits_data;
  wire [1:0]   slave2_r_bits_resp_0 = slave2_r_bits_resp;
  wire         slave2_r_bits_last_0 = slave2_r_bits_last;
  wire         slave3_aw_ready_0 = slave3_aw_ready;
  wire         slave3_w_ready_0 = slave3_w_ready;
  wire         slave3_b_valid_0 = slave3_b_valid;
  wire [7:0]   slave3_b_bits_id_0 = slave3_b_bits_id;
  wire [1:0]   slave3_b_bits_resp_0 = slave3_b_bits_resp;
  wire         slave3_ar_ready_0 = slave3_ar_ready;
  wire         slave3_r_valid_0 = slave3_r_valid;
  wire [7:0]   slave3_r_bits_id_0 = slave3_r_bits_id;
  wire [127:0] slave3_r_bits_data_0 = slave3_r_bits_data;
  wire [1:0]   slave3_r_bits_resp_0 = slave3_r_bits_resp;
  wire         slave3_r_bits_last_0 = slave3_r_bits_last;
  wire         slave4_aw_ready_0 = slave4_aw_ready;
  wire         slave4_w_ready_0 = slave4_w_ready;
  wire         slave4_b_valid_0 = slave4_b_valid;
  wire [7:0]   slave4_b_bits_id_0 = slave4_b_bits_id;
  wire [1:0]   slave4_b_bits_resp_0 = slave4_b_bits_resp;
  wire         slave4_ar_ready_0 = slave4_ar_ready;
  wire         slave4_r_valid_0 = slave4_r_valid;
  wire [7:0]   slave4_r_bits_id_0 = slave4_r_bits_id;
  wire [127:0] slave4_r_bits_data_0 = slave4_r_bits_data;
  wire [1:0]   slave4_r_bits_resp_0 = slave4_r_bits_resp;
  wire         slave4_r_bits_last_0 = slave4_r_bits_last;
  wire         xbar_arFIFOMap_1_0 = 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:111:36
  wire         xbar_arFIFOMap_1_1 = 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:111:36
  wire         xbar_awFIFOMap_1_0 = 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:112:36
  wire         xbar_awFIFOMap_1_1 = 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:112:36
  wire [0:0]   _GEN = '{1'h1};
  wire [7:0]   master1_b_bits_id_0 = 8'h0;
  wire [7:0]   master1_r_bits_id_0 = 8'h0;
  wire         xbar_auto_anon_in_0_b_bits_id = 1'h0;
  wire         xbar_auto_anon_in_0_r_bits_id = 1'h0;
  wire         xbar_anonIn_b_bits_id = 1'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_r_bits_id = 1'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapMasterOut_b_bits_id = 1'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_r_bits_id = 1'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_aw_valid = master1_aw_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   mapMasterOut_aw_bits_len = master1_aw_bits_len_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_aw_bits_size = master1_aw_bits_size_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_aw_bits_burst = master1_aw_bits_burst_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_aw_bits_lock = master1_aw_bits_lock_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_aw_bits_cache = master1_aw_bits_cache_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_aw_bits_prot = master1_aw_bits_prot_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_aw_bits_qos = master1_aw_bits_qos_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_w_valid = master1_w_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] mapMasterOut_w_bits_data = master1_w_bits_data_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [15:0]  mapMasterOut_w_bits_strb = master1_w_bits_strb_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_w_bits_last = master1_w_bits_last_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_b_ready = master1_b_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_ar_valid = master1_ar_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   mapMasterOut_ar_bits_len = master1_ar_bits_len_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_ar_bits_size = master1_ar_bits_size_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_ar_bits_burst = master1_ar_bits_burst_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_ar_bits_lock = master1_ar_bits_lock_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_ar_bits_cache = master1_ar_bits_cache_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_ar_bits_prot = master1_ar_bits_prot_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_ar_bits_qos = master1_ar_bits_qos_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_r_ready = master1_r_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] mapMasterOut_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_aw_valid = master2_aw_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   mapMasterOut_1_aw_bits_len = master2_aw_bits_len_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_1_aw_bits_size = master2_aw_bits_size_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_1_aw_bits_burst = master2_aw_bits_burst_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_aw_bits_lock = master2_aw_bits_lock_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_1_aw_bits_cache = master2_aw_bits_cache_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_1_aw_bits_prot = master2_aw_bits_prot_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_1_aw_bits_qos = master2_aw_bits_qos_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_w_valid = master2_w_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] mapMasterOut_1_w_bits_data = master2_w_bits_data_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [15:0]  mapMasterOut_1_w_bits_strb = master2_w_bits_strb_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_w_bits_last = master2_w_bits_last_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_b_ready = master2_b_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_ar_valid = master2_ar_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   mapMasterOut_1_ar_bits_len = master2_ar_bits_len_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_1_ar_bits_size = master2_ar_bits_size_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_1_ar_bits_burst = master2_ar_bits_burst_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_ar_bits_lock = master2_ar_bits_lock_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_1_ar_bits_cache = master2_ar_bits_cache_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapMasterOut_1_ar_bits_prot = master2_ar_bits_prot_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   mapMasterOut_1_ar_bits_qos = master2_ar_bits_qos_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_r_ready = master2_r_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] mapMasterOut_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   mapMasterOut_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapMasterOut_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         mapSlaveIn_aw_ready = slave1_aw_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_w_ready = slave1_w_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  mapSlaveIn_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_b_valid = slave1_b_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_b_bits_resp = slave1_b_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_ar_ready = slave1_ar_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_r_valid = slave1_r_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_r_bits_data = slave1_r_bits_data_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_r_bits_resp = slave1_r_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_r_bits_last = slave1_r_bits_last_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_aw_ready = slave2_aw_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_w_ready = slave2_w_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  mapSlaveIn_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_b_valid = slave2_b_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_1_b_bits_resp = slave2_b_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_ar_ready = slave2_ar_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_r_valid = slave2_r_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_1_r_bits_data = slave2_r_bits_data_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_1_r_bits_resp = slave2_r_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_1_r_bits_last = slave2_r_bits_last_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_aw_ready = slave3_aw_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_2_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_2_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_2_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_2_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_2_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_2_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_w_ready = slave3_w_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_2_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  mapSlaveIn_2_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_b_valid = slave3_b_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_2_b_bits_resp = slave3_b_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_ar_ready = slave3_ar_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_2_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_2_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_2_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_2_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_2_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_2_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_r_valid = slave3_r_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_2_r_bits_data = slave3_r_bits_data_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_2_r_bits_resp = slave3_r_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_2_r_bits_last = slave3_r_bits_last_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_aw_ready = slave4_aw_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_3_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_3_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_3_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_3_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_3_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_3_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_w_ready = slave4_w_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_3_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  mapSlaveIn_3_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_b_valid = slave4_b_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_3_b_bits_resp = slave4_b_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_ar_ready = slave4_ar_ready_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   mapSlaveIn_3_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_3_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_3_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_3_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   mapSlaveIn_3_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   mapSlaveIn_3_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_r_valid = slave4_r_valid_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] mapSlaveIn_3_r_bits_data = slave4_r_bits_data_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapSlaveIn_3_r_bits_resp = slave4_r_bits_resp_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapSlaveIn_3_r_bits_last = slave4_r_bits_last_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_aw_ready = xbar_auto_anon_in_1_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_1_aw_valid = xbar_auto_anon_in_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapMasterOut_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_anonIn_1_aw_bits_id = xbar_auto_anon_in_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  mapMasterOut_1_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar__requestAWIO_T_20 = xbar_auto_anon_in_1_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_anonIn_1_aw_bits_len = xbar_auto_anon_in_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_1_aw_bits_size = xbar_auto_anon_in_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonIn_1_aw_bits_burst = xbar_auto_anon_in_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_aw_bits_lock = xbar_auto_anon_in_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_1_aw_bits_cache = xbar_auto_anon_in_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_1_aw_bits_prot = xbar_auto_anon_in_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_1_aw_bits_qos = xbar_auto_anon_in_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_w_ready = xbar_auto_anon_in_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_1_w_valid = xbar_auto_anon_in_1_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] xbar_anonIn_1_w_bits_data = xbar_auto_anon_in_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  xbar_anonIn_1_w_bits_strb = xbar_auto_anon_in_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_w_bits_last = xbar_auto_anon_in_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_b_ready = xbar_auto_anon_in_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonIn_1_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_b_valid = xbar_auto_anon_in_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_anonIn_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapMasterOut_1_b_bits_id = xbar_auto_anon_in_1_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_b_bits_resp = xbar_auto_anon_in_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapMasterOut_1_ar_ready = xbar_auto_anon_in_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_1_ar_valid = xbar_auto_anon_in_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapMasterOut_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_anonIn_1_ar_bits_id = xbar_auto_anon_in_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  mapMasterOut_1_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar__requestARIO_T_20 = xbar_auto_anon_in_1_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_anonIn_1_ar_bits_len = xbar_auto_anon_in_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_1_ar_bits_size = xbar_auto_anon_in_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonIn_1_ar_bits_burst = xbar_auto_anon_in_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_ar_bits_lock = xbar_auto_anon_in_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_1_ar_bits_cache = xbar_auto_anon_in_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_1_ar_bits_prot = xbar_auto_anon_in_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_1_ar_bits_qos = xbar_auto_anon_in_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_r_ready = xbar_auto_anon_in_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonIn_1_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_r_valid = xbar_auto_anon_in_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_anonIn_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   mapMasterOut_1_r_bits_id = xbar_auto_anon_in_1_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_anonIn_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_r_bits_data = xbar_auto_anon_in_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_r_bits_resp = xbar_auto_anon_in_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_1_r_bits_last = xbar_auto_anon_in_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapMasterOut_aw_ready = xbar_auto_anon_in_0_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_aw_valid = xbar_auto_anon_in_0_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapMasterOut_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_aw_bits_id = xbar_auto_anon_in_0_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  mapMasterOut_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar__requestAWIO_T = xbar_auto_anon_in_0_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_anonIn_aw_bits_len = xbar_auto_anon_in_0_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_aw_bits_size = xbar_auto_anon_in_0_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonIn_aw_bits_burst = xbar_auto_anon_in_0_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_aw_bits_lock = xbar_auto_anon_in_0_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_aw_bits_cache = xbar_auto_anon_in_0_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_aw_bits_prot = xbar_auto_anon_in_0_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_aw_bits_qos = xbar_auto_anon_in_0_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_w_ready = xbar_auto_anon_in_0_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_w_valid = xbar_auto_anon_in_0_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] xbar_anonIn_w_bits_data = xbar_auto_anon_in_0_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  xbar_anonIn_w_bits_strb = xbar_auto_anon_in_0_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_w_bits_last = xbar_auto_anon_in_0_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_b_ready = xbar_auto_anon_in_0_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_b_valid = xbar_auto_anon_in_0_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_anonIn_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_b_bits_resp = xbar_auto_anon_in_0_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapMasterOut_ar_ready = xbar_auto_anon_in_0_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_ar_valid = xbar_auto_anon_in_0_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         mapMasterOut_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_ar_bits_id = xbar_auto_anon_in_0_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  mapMasterOut_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar__requestARIO_T = xbar_auto_anon_in_0_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_anonIn_ar_bits_len = xbar_auto_anon_in_0_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_ar_bits_size = xbar_auto_anon_in_0_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonIn_ar_bits_burst = xbar_auto_anon_in_0_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_ar_bits_lock = xbar_auto_anon_in_0_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_ar_bits_cache = xbar_auto_anon_in_0_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonIn_ar_bits_prot = xbar_auto_anon_in_0_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonIn_ar_bits_qos = xbar_auto_anon_in_0_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_r_ready = xbar_auto_anon_in_0_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonIn_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_r_valid = xbar_auto_anon_in_0_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_anonIn_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonIn_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_r_bits_data = xbar_auto_anon_in_0_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonIn_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_r_bits_resp = xbar_auto_anon_in_0_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapMasterOut_r_bits_last = xbar_auto_anon_in_0_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_2_aw_ready = xbar_auto_anon_out_3_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_2_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_x1_anonOut_2_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_aw_valid = xbar_auto_anon_out_3_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  xbar_x1_anonOut_2_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_3_aw_bits_id = xbar_auto_anon_out_3_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_x1_anonOut_2_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  mapSlaveIn_3_aw_bits_addr = xbar_auto_anon_out_3_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_2_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_aw_bits_len = xbar_auto_anon_out_3_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_x1_anonOut_2_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_aw_bits_size = xbar_auto_anon_out_3_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_aw_bits_burst = xbar_auto_anon_out_3_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_2_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_aw_bits_lock = xbar_auto_anon_out_3_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_2_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_aw_bits_cache = xbar_auto_anon_out_3_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_2_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_aw_bits_prot = xbar_auto_anon_out_3_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_3_aw_bits_qos = xbar_auto_anon_out_3_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_w_ready = xbar_auto_anon_out_3_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_2_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_x1_anonOut_2_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_w_valid = xbar_auto_anon_out_3_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  xbar_x1_anonOut_2_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_w_bits_data = xbar_auto_anon_out_3_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_w_bits_strb = xbar_auto_anon_out_3_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_w_bits_last = xbar_auto_anon_out_3_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_3_b_ready = xbar_auto_anon_out_3_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_b_valid = xbar_auto_anon_out_3_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_3_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar__requestBOI_uncommonBits_T_3 = xbar_auto_anon_out_3_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_x1_anonOut_2_b_bits_resp = xbar_auto_anon_out_3_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_2_ar_ready = xbar_auto_anon_out_3_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_2_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_x1_anonOut_2_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_valid = xbar_auto_anon_out_3_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  xbar_x1_anonOut_2_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_3_ar_bits_id = xbar_auto_anon_out_3_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_x1_anonOut_2_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  mapSlaveIn_3_ar_bits_addr = xbar_auto_anon_out_3_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_2_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_bits_len = xbar_auto_anon_out_3_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_x1_anonOut_2_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_bits_size = xbar_auto_anon_out_3_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_bits_burst = xbar_auto_anon_out_3_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_2_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_bits_lock = xbar_auto_anon_out_3_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_2_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_bits_cache = xbar_auto_anon_out_3_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_2_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_bits_prot = xbar_auto_anon_out_3_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_3_ar_bits_qos = xbar_auto_anon_out_3_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_3_r_ready = xbar_auto_anon_out_3_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_2_r_valid = xbar_auto_anon_out_3_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_3_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar__requestROI_uncommonBits_T_3 = xbar_auto_anon_out_3_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_x1_anonOut_2_r_bits_data = xbar_auto_anon_out_3_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_x1_anonOut_2_r_bits_resp = xbar_auto_anon_out_3_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_2_r_bits_last = xbar_auto_anon_out_3_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_1_aw_ready = xbar_auto_anon_out_2_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_x1_anonOut_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_aw_valid = xbar_auto_anon_out_2_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  xbar_x1_anonOut_1_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_2_aw_bits_id = xbar_auto_anon_out_2_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_x1_anonOut_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  mapSlaveIn_2_aw_bits_addr = xbar_auto_anon_out_2_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_aw_bits_len = xbar_auto_anon_out_2_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_x1_anonOut_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_aw_bits_size = xbar_auto_anon_out_2_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_aw_bits_burst = xbar_auto_anon_out_2_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_aw_bits_lock = xbar_auto_anon_out_2_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_aw_bits_cache = xbar_auto_anon_out_2_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_aw_bits_prot = xbar_auto_anon_out_2_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_2_aw_bits_qos = xbar_auto_anon_out_2_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_w_ready = xbar_auto_anon_out_2_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_1_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_x1_anonOut_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_w_valid = xbar_auto_anon_out_2_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  xbar_x1_anonOut_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_w_bits_data = xbar_auto_anon_out_2_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_w_bits_strb = xbar_auto_anon_out_2_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_w_bits_last = xbar_auto_anon_out_2_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_2_b_ready = xbar_auto_anon_out_2_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_b_valid = xbar_auto_anon_out_2_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_2_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar__requestBOI_uncommonBits_T_2 = xbar_auto_anon_out_2_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_x1_anonOut_1_b_bits_resp = xbar_auto_anon_out_2_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_1_ar_ready = xbar_auto_anon_out_2_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_x1_anonOut_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_valid = xbar_auto_anon_out_2_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  xbar_x1_anonOut_1_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_2_ar_bits_id = xbar_auto_anon_out_2_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_x1_anonOut_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  mapSlaveIn_2_ar_bits_addr = xbar_auto_anon_out_2_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_bits_len = xbar_auto_anon_out_2_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_x1_anonOut_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_bits_size = xbar_auto_anon_out_2_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_bits_burst = xbar_auto_anon_out_2_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_bits_lock = xbar_auto_anon_out_2_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_bits_cache = xbar_auto_anon_out_2_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_bits_prot = xbar_auto_anon_out_2_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_2_ar_bits_qos = xbar_auto_anon_out_2_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_2_r_ready = xbar_auto_anon_out_2_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_1_r_valid = xbar_auto_anon_out_2_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_2_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar__requestROI_uncommonBits_T_2 = xbar_auto_anon_out_2_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_x1_anonOut_1_r_bits_data = xbar_auto_anon_out_2_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_x1_anonOut_1_r_bits_resp = xbar_auto_anon_out_2_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_1_r_bits_last = xbar_auto_anon_out_2_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_aw_ready = xbar_auto_anon_out_1_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_x1_anonOut_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_aw_valid = xbar_auto_anon_out_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [28:0]  xbar_x1_anonOut_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_1_aw_bits_id = xbar_auto_anon_out_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_x1_anonOut_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [28:0]  mapSlaveIn_1_aw_bits_addr = xbar_auto_anon_out_1_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_aw_bits_len = xbar_auto_anon_out_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_x1_anonOut_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_aw_bits_size = xbar_auto_anon_out_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_aw_bits_burst = xbar_auto_anon_out_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_aw_bits_lock = xbar_auto_anon_out_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_aw_bits_cache = xbar_auto_anon_out_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_aw_bits_prot = xbar_auto_anon_out_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_1_aw_bits_qos = xbar_auto_anon_out_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_w_ready = xbar_auto_anon_out_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_x1_anonOut_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_w_valid = xbar_auto_anon_out_1_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  xbar_x1_anonOut_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_w_bits_data = xbar_auto_anon_out_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_w_bits_strb = xbar_auto_anon_out_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_w_bits_last = xbar_auto_anon_out_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_1_b_ready = xbar_auto_anon_out_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_b_valid = xbar_auto_anon_out_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_1_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_b_bits_id = xbar_auto_anon_out_1_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_x1_anonOut_b_bits_resp = xbar_auto_anon_out_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_ar_ready = xbar_auto_anon_out_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_x1_anonOut_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_valid = xbar_auto_anon_out_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [28:0]  xbar_x1_anonOut_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_1_ar_bits_id = xbar_auto_anon_out_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_x1_anonOut_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [28:0]  mapSlaveIn_1_ar_bits_addr = xbar_auto_anon_out_1_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_bits_len = xbar_auto_anon_out_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_x1_anonOut_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_bits_size = xbar_auto_anon_out_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_bits_burst = xbar_auto_anon_out_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_bits_lock = xbar_auto_anon_out_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_bits_cache = xbar_auto_anon_out_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_x1_anonOut_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_bits_prot = xbar_auto_anon_out_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_1_ar_bits_qos = xbar_auto_anon_out_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_1_r_ready = xbar_auto_anon_out_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_x1_anonOut_r_valid = xbar_auto_anon_out_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_1_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_x1_anonOut_r_bits_id = xbar_auto_anon_out_1_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_x1_anonOut_r_bits_data = xbar_auto_anon_out_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_x1_anonOut_r_bits_resp = xbar_auto_anon_out_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_x1_anonOut_r_bits_last = xbar_auto_anon_out_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonOut_aw_ready = xbar_auto_anon_out_0_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonOut_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_anonOut_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_aw_valid = xbar_auto_anon_out_0_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [27:0]  xbar_anonOut_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_aw_bits_id = xbar_auto_anon_out_0_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_anonOut_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [27:0]  mapSlaveIn_aw_bits_addr = xbar_auto_anon_out_0_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonOut_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_aw_bits_len = xbar_auto_anon_out_0_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonOut_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_aw_bits_size = xbar_auto_anon_out_0_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_aw_bits_burst = xbar_auto_anon_out_0_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonOut_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_aw_bits_lock = xbar_auto_anon_out_0_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonOut_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_aw_bits_cache = xbar_auto_anon_out_0_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonOut_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_aw_bits_prot = xbar_auto_anon_out_0_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_aw_bits_qos = xbar_auto_anon_out_0_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_w_ready = xbar_auto_anon_out_0_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonOut_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_anonOut_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_w_valid = xbar_auto_anon_out_0_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  xbar_anonOut_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_w_bits_data = xbar_auto_anon_out_0_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_w_bits_strb = xbar_auto_anon_out_0_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_w_bits_last = xbar_auto_anon_out_0_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_b_ready = xbar_auto_anon_out_0_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_b_valid = xbar_auto_anon_out_0_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonOut_b_bits_id = xbar_auto_anon_out_0_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_anonOut_b_bits_resp = xbar_auto_anon_out_0_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonOut_ar_ready = xbar_auto_anon_out_0_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonOut_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_anonOut_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_valid = xbar_auto_anon_out_0_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [27:0]  xbar_anonOut_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_ar_bits_id = xbar_auto_anon_out_0_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   xbar_anonOut_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [27:0]  mapSlaveIn_ar_bits_addr = xbar_auto_anon_out_0_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonOut_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_bits_len = xbar_auto_anon_out_0_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_anonOut_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_bits_size = xbar_auto_anon_out_0_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_bits_burst = xbar_auto_anon_out_0_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonOut_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_bits_lock = xbar_auto_anon_out_0_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonOut_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_bits_cache = xbar_auto_anon_out_0_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   xbar_anonOut_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_bits_prot = xbar_auto_anon_out_0_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign mapSlaveIn_ar_bits_qos = xbar_auto_anon_out_0_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapSlaveIn_r_ready = xbar_auto_anon_out_0_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_anonOut_r_valid = xbar_auto_anon_out_0_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   mapSlaveIn_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   xbar_anonOut_r_bits_id = xbar_auto_anon_out_0_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_anonOut_r_bits_data = xbar_auto_anon_out_0_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_anonOut_r_bits_resp = xbar_auto_anon_out_0_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_anonOut_r_bits_last = xbar_auto_anon_out_0_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_ready = xbar_anonIn_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  xbar_in_0_aw_bits_addr = xbar__requestAWIO_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [7:0]   xbar_in_0_aw_bits_len = xbar_anonIn_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_0_aw_bits_size = xbar_anonIn_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [1:0]   xbar_in_0_aw_bits_burst = xbar_anonIn_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_aw_bits_lock = xbar_anonIn_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_0_aw_bits_cache = xbar_anonIn_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_0_aw_bits_prot = xbar_anonIn_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_0_aw_bits_qos = xbar_anonIn_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_0_w_ready = xbar_anonIn_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] xbar_in_0_w_bits_data = xbar_anonIn_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [15:0]  xbar_in_0_w_bits_strb = xbar_anonIn_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_w_bits_last = xbar_anonIn_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_b_ready = xbar_anonIn_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_b_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_0_b_valid = xbar_anonIn_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_in_0_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_0_b_bits_resp = xbar_anonIn_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_in_0_ar_ready = xbar_anonIn_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [29:0]  xbar_in_0_ar_bits_addr = xbar__requestARIO_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [7:0]   xbar_in_0_ar_bits_len = xbar_anonIn_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_0_ar_bits_size = xbar_anonIn_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [1:0]   xbar_in_0_ar_bits_burst = xbar_anonIn_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_ar_bits_lock = xbar_anonIn_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_0_ar_bits_cache = xbar_anonIn_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_0_ar_bits_prot = xbar_anonIn_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_0_ar_bits_qos = xbar_anonIn_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_r_ready = xbar_anonIn_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_r_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_0_r_valid = xbar_anonIn_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] xbar_in_0_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_0_r_bits_data = xbar_anonIn_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_in_0_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_0_r_bits_resp = xbar_anonIn_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_in_0_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_0_r_bits_last = xbar_anonIn_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_in_1_aw_ready = xbar_anonIn_1_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_awSel_shiftAmount = xbar_anonIn_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/chisel3/util/OneHot.scala:64:49
  wire [29:0]  xbar_in_1_aw_bits_addr = xbar__requestAWIO_T_20;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [7:0]   xbar_in_1_aw_bits_len = xbar_anonIn_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_1_aw_bits_size = xbar_anonIn_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [1:0]   xbar_in_1_aw_bits_burst = xbar_anonIn_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_aw_bits_lock = xbar_anonIn_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_1_aw_bits_cache = xbar_anonIn_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_1_aw_bits_prot = xbar_anonIn_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_1_aw_bits_qos = xbar_anonIn_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_1_w_ready = xbar_anonIn_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] xbar_in_1_w_bits_data = xbar_anonIn_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [15:0]  xbar_in_1_w_bits_strb = xbar_anonIn_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_w_bits_last = xbar_anonIn_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_b_ready = xbar_anonIn_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_b_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_1_b_valid = xbar_anonIn_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_in_1_b_bits_id = xbar_anonIn_1_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_in_1_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [1:0]   xbar_bSel_shiftAmount = xbar_anonIn_1_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/chisel3/util/OneHot.scala:64:49
  assign xbar_auto_anon_in_1_b_bits_resp = xbar_anonIn_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_in_1_ar_ready = xbar_anonIn_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_arSel_shiftAmount = xbar_anonIn_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/chisel3/util/OneHot.scala:64:49
  wire [29:0]  xbar_in_1_ar_bits_addr = xbar__requestARIO_T_20;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [7:0]   xbar_in_1_ar_bits_len = xbar_anonIn_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_1_ar_bits_size = xbar_anonIn_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [1:0]   xbar_in_1_ar_bits_burst = xbar_anonIn_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_ar_bits_lock = xbar_anonIn_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_1_ar_bits_cache = xbar_anonIn_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_in_1_ar_bits_prot = xbar_anonIn_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [3:0]   xbar_in_1_ar_bits_qos = xbar_anonIn_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_r_ready = xbar_anonIn_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_r_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_1_r_valid = xbar_anonIn_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_in_1_r_bits_id = xbar_anonIn_1_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] xbar_in_1_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [1:0]   xbar_rSel_shiftAmount = xbar_anonIn_1_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/chisel3/util/OneHot.scala:64:49
  assign xbar_auto_anon_in_1_r_bits_data = xbar_anonIn_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   xbar_in_1_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_1_r_bits_resp = xbar_anonIn_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         xbar_in_1_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_auto_anon_in_1_r_bits_last = xbar_anonIn_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_aw_valid = xbar_anonOut_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_0_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_id = xbar_anonOut_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_0_aw_bits_addr = xbar_anonOut_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_0_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_len = xbar_anonOut_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_0_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_size = xbar_anonOut_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_0_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_burst = xbar_anonOut_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_0_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_lock = xbar_anonOut_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_0_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_cache = xbar_anonOut_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_0_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_prot = xbar_anonOut_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_0_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_aw_bits_qos = xbar_anonOut_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_0_w_valid = xbar_anonOut_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_out_0_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_w_bits_data = xbar_anonOut_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [15:0]  xbar_out_0_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_w_bits_strb = xbar_anonOut_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_0_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_w_bits_last = xbar_anonOut_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_0_b_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_b_ready = xbar_anonOut_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_0_b_valid = xbar_anonOut_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_0_b_bits_id = xbar_anonOut_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_0_b_bits_resp = xbar_anonOut_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_0_ar_ready = xbar_anonOut_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_0_ar_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_valid = xbar_anonOut_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_0_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_id = xbar_anonOut_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_0_ar_bits_addr = xbar_anonOut_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_0_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_len = xbar_anonOut_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_0_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_size = xbar_anonOut_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_0_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_burst = xbar_anonOut_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_0_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_lock = xbar_anonOut_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_0_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_cache = xbar_anonOut_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_0_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_prot = xbar_anonOut_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_0_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_ar_bits_qos = xbar_anonOut_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_0_r_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_0_r_ready = xbar_anonOut_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_0_r_valid = xbar_anonOut_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_0_r_bits_id = xbar_anonOut_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [127:0] xbar_out_0_r_bits_data = xbar_anonOut_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_0_r_bits_resp = xbar_anonOut_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_0_r_bits_last = xbar_anonOut_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_valid = xbar_x1_anonOut_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_1_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_id = xbar_x1_anonOut_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_1_aw_bits_addr = xbar_x1_anonOut_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_1_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_len = xbar_x1_anonOut_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_1_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_size = xbar_x1_anonOut_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_1_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_burst = xbar_x1_anonOut_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_1_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_lock = xbar_x1_anonOut_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_1_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_cache = xbar_x1_anonOut_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_1_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_prot = xbar_x1_anonOut_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_1_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_aw_bits_qos = xbar_x1_anonOut_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_1_w_valid = xbar_x1_anonOut_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_out_1_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_w_bits_data = xbar_x1_anonOut_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [15:0]  xbar_out_1_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_w_bits_strb = xbar_x1_anonOut_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_1_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_w_bits_last = xbar_x1_anonOut_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_1_b_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_b_ready = xbar_x1_anonOut_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_1_b_valid = xbar_x1_anonOut_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_1_b_bits_id = xbar_x1_anonOut_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_1_b_bits_resp = xbar_x1_anonOut_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_1_ar_ready = xbar_x1_anonOut_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_1_ar_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_valid = xbar_x1_anonOut_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_1_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_id = xbar_x1_anonOut_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_1_ar_bits_addr = xbar_x1_anonOut_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_1_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_len = xbar_x1_anonOut_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_1_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_size = xbar_x1_anonOut_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_1_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_burst = xbar_x1_anonOut_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_1_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_lock = xbar_x1_anonOut_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_1_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_cache = xbar_x1_anonOut_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_1_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_prot = xbar_x1_anonOut_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_1_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_ar_bits_qos = xbar_x1_anonOut_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_1_r_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_1_r_ready = xbar_x1_anonOut_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_1_r_valid = xbar_x1_anonOut_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_1_r_bits_id = xbar_x1_anonOut_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [127:0] xbar_out_1_r_bits_data = xbar_x1_anonOut_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_1_r_bits_resp = xbar_x1_anonOut_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_1_r_bits_last = xbar_x1_anonOut_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_valid = xbar_x1_anonOut_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_2_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_id = xbar_x1_anonOut_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar_out_2_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_addr = xbar_x1_anonOut_1_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_2_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_len = xbar_x1_anonOut_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_2_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_size = xbar_x1_anonOut_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_2_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_burst = xbar_x1_anonOut_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_2_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_lock = xbar_x1_anonOut_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_2_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_cache = xbar_x1_anonOut_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_2_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_prot = xbar_x1_anonOut_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_2_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_aw_bits_qos = xbar_x1_anonOut_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_2_w_valid = xbar_x1_anonOut_1_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_out_2_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_w_bits_data = xbar_x1_anonOut_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [15:0]  xbar_out_2_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_w_bits_strb = xbar_x1_anonOut_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_2_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_w_bits_last = xbar_x1_anonOut_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_2_b_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_b_ready = xbar_x1_anonOut_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_2_b_valid = xbar_x1_anonOut_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_2_b_bits_id = xbar__requestBOI_uncommonBits_T_2;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_2_b_bits_resp = xbar_x1_anonOut_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_2_ar_ready = xbar_x1_anonOut_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_2_ar_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_valid = xbar_x1_anonOut_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_2_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_id = xbar_x1_anonOut_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar_out_2_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_addr = xbar_x1_anonOut_1_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_2_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_len = xbar_x1_anonOut_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_2_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_size = xbar_x1_anonOut_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_2_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_burst = xbar_x1_anonOut_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_2_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_lock = xbar_x1_anonOut_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_2_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_cache = xbar_x1_anonOut_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_2_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_prot = xbar_x1_anonOut_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_2_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_ar_bits_qos = xbar_x1_anonOut_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_2_r_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_2_r_ready = xbar_x1_anonOut_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_2_r_valid = xbar_x1_anonOut_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_2_r_bits_id = xbar__requestROI_uncommonBits_T_2;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [127:0] xbar_out_2_r_bits_data = xbar_x1_anonOut_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_2_r_bits_resp = xbar_x1_anonOut_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_2_r_bits_last = xbar_x1_anonOut_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_valid = xbar_x1_anonOut_2_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_3_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_id = xbar_x1_anonOut_2_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar_out_3_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_addr = xbar_x1_anonOut_2_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_3_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_len = xbar_x1_anonOut_2_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_3_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_size = xbar_x1_anonOut_2_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_3_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_burst = xbar_x1_anonOut_2_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_3_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_lock = xbar_x1_anonOut_2_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_3_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_cache = xbar_x1_anonOut_2_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_3_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_prot = xbar_x1_anonOut_2_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_3_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_aw_bits_qos = xbar_x1_anonOut_2_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_3_w_valid = xbar_x1_anonOut_2_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] xbar_out_3_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_w_bits_data = xbar_x1_anonOut_2_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [15:0]  xbar_out_3_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_w_bits_strb = xbar_x1_anonOut_2_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_3_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_w_bits_last = xbar_x1_anonOut_2_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_3_b_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_b_ready = xbar_x1_anonOut_2_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_3_b_valid = xbar_x1_anonOut_2_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_3_b_bits_id = xbar__requestBOI_uncommonBits_T_3;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_3_b_bits_resp = xbar_x1_anonOut_2_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_3_ar_ready = xbar_x1_anonOut_2_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_3_ar_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_valid = xbar_x1_anonOut_2_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_3_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_id = xbar_x1_anonOut_2_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [29:0]  xbar_out_3_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_addr = xbar_x1_anonOut_2_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [7:0]   xbar_out_3_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_len = xbar_x1_anonOut_2_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_3_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_size = xbar_x1_anonOut_2_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   xbar_out_3_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_burst = xbar_x1_anonOut_2_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_3_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_lock = xbar_x1_anonOut_2_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_3_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_cache = xbar_x1_anonOut_2_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [2:0]   xbar_out_3_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_prot = xbar_x1_anonOut_2_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [3:0]   xbar_out_3_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_ar_bits_qos = xbar_x1_anonOut_2_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_3_r_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_auto_anon_out_3_r_ready = xbar_x1_anonOut_2_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         xbar_out_3_r_valid = xbar_x1_anonOut_2_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_out_3_r_bits_id = xbar__requestROI_uncommonBits_T_3;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [127:0] xbar_out_3_r_bits_data = xbar_x1_anonOut_2_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [1:0]   xbar_out_3_r_bits_resp = xbar_x1_anonOut_2_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_out_3_r_bits_last = xbar_x1_anonOut_2_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  reg          xbar_awIn_0_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awIn_0_wrap = xbar_awIn_0_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awIn_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awIn_0_wrap_1 = xbar_awIn_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awIn_0_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
  wire         xbar_awIn_0_ptr_match =
    xbar_awIn_0_enq_ptr_value == xbar_awIn_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:261:33
  wire         xbar_awIn_0_empty = xbar_awIn_0_ptr_match & ~xbar_awIn_0_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :262:{25,28}
  wire         xbar_awIn_0_full = xbar_awIn_0_ptr_match & xbar_awIn_0_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :263:24
  wire         xbar_awIn_0_io_enq_ready = ~xbar_awIn_0_full;	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :287:19
  wire         xbar_awIn_0_io_enq_valid;
  wire [3:0]   xbar_awIn_0_io_enq_bits;
  wire         xbar_awIn_0_io_deq_valid = xbar_awIn_0_io_enq_valid | ~xbar_awIn_0_empty;	// src/main/scala/chisel3/util/Decoupled.scala:262:25, :286:{16,19}, :298:{24,39}
  wire [3:0]   xbar_awIn_0_io_deq_bits =
    xbar_awIn_0_empty ? xbar_awIn_0_io_enq_bits : _ram_ext_R0_data_4;	// src/main/scala/chisel3/util/Decoupled.scala:257:91, :262:25, :294:17, :299:17, :300:19
  wire         xbar_awIn_0_io_deq_ready;
  wire         xbar_awIn_0_do_deq =
    ~xbar_awIn_0_empty & xbar_awIn_0_io_deq_ready & xbar_awIn_0_io_deq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :265:27, :299:17, :301:14
  wire         xbar_awIn_0_do_enq =
    ~(xbar_awIn_0_empty & xbar_awIn_0_io_deq_ready) & xbar_awIn_0_io_enq_ready
    & xbar_awIn_0_io_enq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :264:27, :299:17, :302:{26,35}
  wire         xbar_awIn_0_ptr_diff =
    xbar_awIn_0_enq_ptr_value - xbar_awIn_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:310:32
  wire [1:0]   xbar_awIn_0_io_count = {xbar_awIn_0_full, xbar_awIn_0_ptr_diff};	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :310:32, :313:62
  reg          xbar_awIn_1_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awIn_1_wrap = xbar_awIn_1_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awIn_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awIn_1_wrap_1 = xbar_awIn_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awIn_1_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
  wire         xbar_awIn_1_ptr_match =
    xbar_awIn_1_enq_ptr_value == xbar_awIn_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:261:33
  wire         xbar_awIn_1_empty = xbar_awIn_1_ptr_match & ~xbar_awIn_1_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :262:{25,28}
  wire         xbar_awIn_1_full = xbar_awIn_1_ptr_match & xbar_awIn_1_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :263:24
  wire         xbar_awIn_1_io_enq_ready = ~xbar_awIn_1_full;	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :287:19
  wire         xbar_awIn_1_io_enq_valid;
  wire [3:0]   xbar_awIn_1_io_enq_bits;
  wire         xbar_awIn_1_io_deq_valid = xbar_awIn_1_io_enq_valid | ~xbar_awIn_1_empty;	// src/main/scala/chisel3/util/Decoupled.scala:262:25, :286:{16,19}, :298:{24,39}
  wire [3:0]   xbar_awIn_1_io_deq_bits =
    xbar_awIn_1_empty ? xbar_awIn_1_io_enq_bits : _ram_ext_R0_data_3;	// src/main/scala/chisel3/util/Decoupled.scala:257:91, :262:25, :294:17, :299:17, :300:19
  wire         xbar_awIn_1_io_deq_ready;
  wire         xbar_awIn_1_do_deq =
    ~xbar_awIn_1_empty & xbar_awIn_1_io_deq_ready & xbar_awIn_1_io_deq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :265:27, :299:17, :301:14
  wire         xbar_awIn_1_do_enq =
    ~(xbar_awIn_1_empty & xbar_awIn_1_io_deq_ready) & xbar_awIn_1_io_enq_ready
    & xbar_awIn_1_io_enq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :264:27, :299:17, :302:{26,35}
  wire         xbar_awIn_1_ptr_diff =
    xbar_awIn_1_enq_ptr_value - xbar_awIn_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:310:32
  wire [1:0]   xbar_awIn_1_io_count = {xbar_awIn_1_full, xbar_awIn_1_ptr_diff};	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :310:32, :313:62
  reg          xbar_awOut_0_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_0_wrap = xbar_awOut_0_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_0_wrap_1 = xbar_awOut_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_0_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
  wire         xbar_awOut_0_ptr_match =
    xbar_awOut_0_enq_ptr_value == xbar_awOut_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:261:33
  wire         xbar_awOut_0_empty = xbar_awOut_0_ptr_match & ~xbar_awOut_0_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :262:{25,28}
  wire         xbar_awOut_0_full = xbar_awOut_0_ptr_match & xbar_awOut_0_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :263:24
  wire         xbar_awOut_0_io_enq_ready = ~xbar_awOut_0_full;	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :287:19
  wire         xbar_awOut_0_io_enq_valid;
  wire [1:0]   xbar_awOut_0_io_enq_bits;
  wire         xbar_awOut_0_io_deq_valid =
    xbar_awOut_0_io_enq_valid | ~xbar_awOut_0_empty;	// src/main/scala/chisel3/util/Decoupled.scala:262:25, :286:{16,19}, :298:{24,39}
  wire [1:0]   xbar_awOut_0_io_deq_bits =
    xbar_awOut_0_empty ? xbar_awOut_0_io_enq_bits : _ram_ext_R0_data_2;	// src/main/scala/chisel3/util/Decoupled.scala:257:91, :262:25, :294:17, :299:17, :300:19
  wire         xbar_awOut_0_io_deq_ready;
  wire         xbar_awOut_0_do_deq =
    ~xbar_awOut_0_empty & xbar_awOut_0_io_deq_ready & xbar_awOut_0_io_deq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :265:27, :299:17, :301:14
  wire         xbar_awOut_0_do_enq =
    ~(xbar_awOut_0_empty & xbar_awOut_0_io_deq_ready) & xbar_awOut_0_io_enq_ready
    & xbar_awOut_0_io_enq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :264:27, :299:17, :302:{26,35}
  wire         xbar_awOut_0_ptr_diff =
    xbar_awOut_0_enq_ptr_value - xbar_awOut_0_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:310:32
  wire [1:0]   xbar_awOut_0_io_count = {xbar_awOut_0_full, xbar_awOut_0_ptr_diff};	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :310:32, :313:62
  reg          xbar_awOut_1_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_1_wrap = xbar_awOut_1_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_1_wrap_1 = xbar_awOut_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_1_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
  wire         xbar_awOut_1_ptr_match =
    xbar_awOut_1_enq_ptr_value == xbar_awOut_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:261:33
  wire         xbar_awOut_1_empty = xbar_awOut_1_ptr_match & ~xbar_awOut_1_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :262:{25,28}
  wire         xbar_awOut_1_full = xbar_awOut_1_ptr_match & xbar_awOut_1_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :263:24
  wire         xbar_awOut_1_io_enq_ready = ~xbar_awOut_1_full;	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :287:19
  wire         xbar_awOut_1_io_enq_valid;
  wire [1:0]   xbar_awOut_1_io_enq_bits;
  wire         xbar_awOut_1_io_deq_valid =
    xbar_awOut_1_io_enq_valid | ~xbar_awOut_1_empty;	// src/main/scala/chisel3/util/Decoupled.scala:262:25, :286:{16,19}, :298:{24,39}
  wire [1:0]   xbar_awOut_1_io_deq_bits =
    xbar_awOut_1_empty ? xbar_awOut_1_io_enq_bits : _ram_ext_R0_data_1;	// src/main/scala/chisel3/util/Decoupled.scala:257:91, :262:25, :294:17, :299:17, :300:19
  wire         xbar_awOut_1_io_deq_ready;
  wire         xbar_awOut_1_do_deq =
    ~xbar_awOut_1_empty & xbar_awOut_1_io_deq_ready & xbar_awOut_1_io_deq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :265:27, :299:17, :301:14
  wire         xbar_awOut_1_do_enq =
    ~(xbar_awOut_1_empty & xbar_awOut_1_io_deq_ready) & xbar_awOut_1_io_enq_ready
    & xbar_awOut_1_io_enq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :264:27, :299:17, :302:{26,35}
  wire         xbar_awOut_1_ptr_diff =
    xbar_awOut_1_enq_ptr_value - xbar_awOut_1_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:310:32
  wire [1:0]   xbar_awOut_1_io_count = {xbar_awOut_1_full, xbar_awOut_1_ptr_diff};	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :310:32, :313:62
  reg          xbar_awOut_2_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_2_wrap = xbar_awOut_2_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_2_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_2_wrap_1 = xbar_awOut_2_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_2_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
  wire         xbar_awOut_2_ptr_match =
    xbar_awOut_2_enq_ptr_value == xbar_awOut_2_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:261:33
  wire         xbar_awOut_2_empty = xbar_awOut_2_ptr_match & ~xbar_awOut_2_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :262:{25,28}
  wire         xbar_awOut_2_full = xbar_awOut_2_ptr_match & xbar_awOut_2_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :263:24
  wire         xbar_awOut_2_io_enq_ready = ~xbar_awOut_2_full;	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :287:19
  wire         xbar_awOut_2_io_enq_valid;
  wire [1:0]   xbar_awOut_2_io_enq_bits;
  wire         xbar_awOut_2_io_deq_valid =
    xbar_awOut_2_io_enq_valid | ~xbar_awOut_2_empty;	// src/main/scala/chisel3/util/Decoupled.scala:262:25, :286:{16,19}, :298:{24,39}
  wire [1:0]   xbar_awOut_2_io_deq_bits =
    xbar_awOut_2_empty ? xbar_awOut_2_io_enq_bits : _ram_ext_R0_data_0;	// src/main/scala/chisel3/util/Decoupled.scala:257:91, :262:25, :294:17, :299:17, :300:19
  wire         xbar_awOut_2_io_deq_ready;
  wire         xbar_awOut_2_do_deq =
    ~xbar_awOut_2_empty & xbar_awOut_2_io_deq_ready & xbar_awOut_2_io_deq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :265:27, :299:17, :301:14
  wire         xbar_awOut_2_do_enq =
    ~(xbar_awOut_2_empty & xbar_awOut_2_io_deq_ready) & xbar_awOut_2_io_enq_ready
    & xbar_awOut_2_io_enq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :264:27, :299:17, :302:{26,35}
  wire         xbar_awOut_2_ptr_diff =
    xbar_awOut_2_enq_ptr_value - xbar_awOut_2_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:310:32
  wire [1:0]   xbar_awOut_2_io_count = {xbar_awOut_2_full, xbar_awOut_2_ptr_diff};	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :310:32, :313:62
  reg          xbar_awOut_3_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_3_wrap = xbar_awOut_3_enq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_3_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40
  wire         xbar_awOut_3_wrap_1 = xbar_awOut_3_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, :73:24
  reg          xbar_awOut_3_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
  wire         xbar_awOut_3_ptr_match =
    xbar_awOut_3_enq_ptr_value == xbar_awOut_3_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:261:33
  wire         xbar_awOut_3_empty = xbar_awOut_3_ptr_match & ~xbar_awOut_3_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :262:{25,28}
  wire         xbar_awOut_3_full = xbar_awOut_3_ptr_match & xbar_awOut_3_maybe_full;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :261:33, :263:24
  wire         xbar_awOut_3_io_enq_ready = ~xbar_awOut_3_full;	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :287:19
  wire         xbar_awOut_3_io_enq_valid;
  wire [1:0]   xbar_awOut_3_io_enq_bits;
  wire         xbar_awOut_3_io_deq_valid =
    xbar_awOut_3_io_enq_valid | ~xbar_awOut_3_empty;	// src/main/scala/chisel3/util/Decoupled.scala:262:25, :286:{16,19}, :298:{24,39}
  wire [1:0]   xbar_awOut_3_io_deq_bits =
    xbar_awOut_3_empty ? xbar_awOut_3_io_enq_bits : _ram_ext_R0_data;	// src/main/scala/chisel3/util/Decoupled.scala:257:91, :262:25, :294:17, :299:17, :300:19
  wire         xbar_awOut_3_io_deq_ready;
  wire         xbar_awOut_3_do_deq =
    ~xbar_awOut_3_empty & xbar_awOut_3_io_deq_ready & xbar_awOut_3_io_deq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :265:27, :299:17, :301:14
  wire         xbar_awOut_3_do_enq =
    ~(xbar_awOut_3_empty & xbar_awOut_3_io_deq_ready) & xbar_awOut_3_io_enq_ready
    & xbar_awOut_3_io_enq_valid;	// src/main/scala/chisel3/util/Decoupled.scala:52:35, :262:25, :264:27, :299:17, :302:{26,35}
  wire         xbar_awOut_3_ptr_diff =
    xbar_awOut_3_enq_ptr_value - xbar_awOut_3_deq_ptr_value;	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:310:32
  wire [1:0]   xbar_awOut_3_io_count = {xbar_awOut_3_full, xbar_awOut_3_ptr_diff};	// src/main/scala/chisel3/util/Decoupled.scala:263:24, :310:32, :313:62
  wire         xbar_requestARIO_0_0 = xbar__requestARIO_T[29:28] == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestARIO_0_1 =
    {xbar__requestARIO_T[29], ~(xbar__requestARIO_T[28])} == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{31,41,46,59}
  wire         xbar_requestARIO_0_2 = xbar__requestARIO_T[29:28] == 2'h2;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestARIO_0_3 = &(xbar__requestARIO_T[29:28]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestARIO_1_0 = xbar__requestARIO_T_20[29:28] == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestARIO_1_1 =
    {xbar__requestARIO_T_20[29], ~(xbar__requestARIO_T_20[28])} == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{31,41,46,59}
  wire         xbar_requestARIO_1_2 = xbar__requestARIO_T_20[29:28] == 2'h2;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestARIO_1_3 = &(xbar__requestARIO_T_20[29:28]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:77:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestAWIO_0_0 = xbar__requestAWIO_T[29:28] == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestAWIO_0_1 =
    {xbar__requestAWIO_T[29], ~(xbar__requestAWIO_T[28])} == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{31,41,46,59}
  wire         xbar_requestAWIO_0_2 = xbar__requestAWIO_T[29:28] == 2'h2;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestAWIO_0_3 = &(xbar__requestAWIO_T[29:28]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestAWIO_1_0 = xbar__requestAWIO_T_20[29:28] == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestAWIO_1_1 =
    {xbar__requestAWIO_T_20[29], ~(xbar__requestAWIO_T_20[28])} == 2'h0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{31,41,46,59}
  wire         xbar_requestAWIO_1_2 = xbar__requestAWIO_T_20[29:28] == 2'h2;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestAWIO_1_3 = &(xbar__requestAWIO_T_20[29:28]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:78:48, src/main/scala/diplomacy/Parameters.scala:137:{41,46,59}
  wire         xbar_requestROI_0_0 = xbar_anonOut_r_bits_id == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestROI_uncommonBits = xbar_anonOut_r_bits_id[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestROI_0_1 = ~(xbar_anonOut_r_bits_id[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire         xbar_requestROI_1_0 = xbar_x1_anonOut_r_bits_id == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestROI_uncommonBits_1 = xbar_x1_anonOut_r_bits_id[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestROI_1_1 = ~(xbar_x1_anonOut_r_bits_id[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire         xbar_requestROI_2_0 = xbar__requestROI_uncommonBits_T_2 == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestROI_uncommonBits_2 = xbar__requestROI_uncommonBits_T_2[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestROI_2_1 = ~(xbar__requestROI_uncommonBits_T_2[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire         xbar_requestROI_3_0 = xbar__requestROI_uncommonBits_T_3 == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestROI_uncommonBits_3 = xbar__requestROI_uncommonBits_T_3[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestROI_3_1 = ~(xbar__requestROI_uncommonBits_T_3[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire         xbar_requestBOI_0_0 = xbar_anonOut_b_bits_id == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestBOI_uncommonBits = xbar_anonOut_b_bits_id[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestBOI_0_1 = ~(xbar_anonOut_b_bits_id[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire         xbar_requestBOI_1_0 = xbar_x1_anonOut_b_bits_id == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestBOI_uncommonBits_1 = xbar_x1_anonOut_b_bits_id[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestBOI_1_1 = ~(xbar_x1_anonOut_b_bits_id[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire         xbar_requestBOI_2_0 = xbar__requestBOI_uncommonBits_T_2 == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestBOI_uncommonBits_2 = xbar__requestBOI_uncommonBits_T_2[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestBOI_2_1 = ~(xbar__requestBOI_uncommonBits_T_2[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire         xbar_requestBOI_3_0 = xbar__requestBOI_uncommonBits_T_3 == 3'h4;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:46:9
  wire [1:0]   xbar_requestBOI_uncommonBits_3 = xbar__requestBOI_uncommonBits_T_3[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:52:56
  wire         xbar_requestBOI_3_1 = ~(xbar__requestBOI_uncommonBits_T_3[2]);	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/diplomacy/Parameters.scala:54:{10,32}, :56:48
  wire [1:0]   _GEN_0 = {xbar_requestAWIO_0_1, xbar_requestAWIO_0_0};	// src/main/scala/amba/axi4/Xbar.scala:78:48, :83:75
  wire [1:0]   xbar_awIn_0_io_enq_bits_lo;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  assign xbar_awIn_0_io_enq_bits_lo = _GEN_0;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  wire [1:0]   xbar_awTag_lo;	// src/main/scala/amba/axi4/Xbar.scala:118:45
  assign xbar_awTag_lo = _GEN_0;	// src/main/scala/amba/axi4/Xbar.scala:83:75, :118:45
  wire [1:0]   _GEN_1 = {xbar_requestAWIO_0_3, xbar_requestAWIO_0_2};	// src/main/scala/amba/axi4/Xbar.scala:78:48, :83:75
  wire [1:0]   xbar_awIn_0_io_enq_bits_hi;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  assign xbar_awIn_0_io_enq_bits_hi = _GEN_1;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  wire [1:0]   xbar_awTag_hi;	// src/main/scala/amba/axi4/Xbar.scala:118:45
  assign xbar_awTag_hi = _GEN_1;	// src/main/scala/amba/axi4/Xbar.scala:83:75, :118:45
  assign xbar_awIn_0_io_enq_bits =
    {xbar_awIn_0_io_enq_bits_hi, xbar_awIn_0_io_enq_bits_lo};	// src/main/scala/amba/axi4/Xbar.scala:83:75
  wire [1:0]   _GEN_2 = {xbar_requestAWIO_1_1, xbar_requestAWIO_1_0};	// src/main/scala/amba/axi4/Xbar.scala:78:48, :83:75
  wire [1:0]   xbar_awIn_1_io_enq_bits_lo;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  assign xbar_awIn_1_io_enq_bits_lo = _GEN_2;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  wire [1:0]   xbar_awTag_lo_2;	// src/main/scala/amba/axi4/Xbar.scala:118:45
  assign xbar_awTag_lo_2 = _GEN_2;	// src/main/scala/amba/axi4/Xbar.scala:83:75, :118:45
  wire [1:0]   _GEN_3 = {xbar_requestAWIO_1_3, xbar_requestAWIO_1_2};	// src/main/scala/amba/axi4/Xbar.scala:78:48, :83:75
  wire [1:0]   xbar_awIn_1_io_enq_bits_hi;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  assign xbar_awIn_1_io_enq_bits_hi = _GEN_3;	// src/main/scala/amba/axi4/Xbar.scala:83:75
  wire [1:0]   xbar_awTag_hi_2;	// src/main/scala/amba/axi4/Xbar.scala:118:45
  assign xbar_awTag_hi_2 = _GEN_3;	// src/main/scala/amba/axi4/Xbar.scala:83:75, :118:45
  assign xbar_awIn_1_io_enq_bits =
    {xbar_awIn_1_io_enq_bits_hi, xbar_awIn_1_io_enq_bits_lo};	// src/main/scala/amba/axi4/Xbar.scala:83:75
  wire         xbar_requestWIO_0_0 = xbar_awIn_0_io_deq_bits[0];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire         xbar_requestWIO_0_1 = xbar_awIn_0_io_deq_bits[1];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire         xbar_requestWIO_0_2 = xbar_awIn_0_io_deq_bits[2];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire         xbar_requestWIO_0_3 = xbar_awIn_0_io_deq_bits[3];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire         xbar_requestWIO_1_0 = xbar_awIn_1_io_deq_bits[0];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire         xbar_requestWIO_1_1 = xbar_awIn_1_io_deq_bits[1];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire         xbar_requestWIO_1_2 = xbar_awIn_1_io_deq_bits[2];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire         xbar_requestWIO_1_3 = xbar_awIn_1_io_deq_bits[3];	// src/main/scala/amba/axi4/Xbar.scala:84:73
  wire [2:0]   xbar_portsAWOI_filtered_0_bits_id = xbar_in_0_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_bits_id = xbar_in_0_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_2_bits_id = xbar_in_0_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_3_bits_id = xbar_in_0_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_0_bits_addr = xbar_in_0_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_1_bits_addr = xbar_in_0_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_2_bits_addr = xbar_in_0_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_3_bits_addr = xbar_in_0_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_0_bits_len = xbar_in_0_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_1_bits_len = xbar_in_0_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_2_bits_len = xbar_in_0_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_3_bits_len = xbar_in_0_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_0_bits_size = xbar_in_0_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_bits_size = xbar_in_0_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_2_bits_size = xbar_in_0_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_3_bits_size = xbar_in_0_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_0_bits_burst = xbar_in_0_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_1_bits_burst = xbar_in_0_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_2_bits_burst = xbar_in_0_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_3_bits_burst = xbar_in_0_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_0_bits_lock = xbar_in_0_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_1_bits_lock = xbar_in_0_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_2_bits_lock = xbar_in_0_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_3_bits_lock = xbar_in_0_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_0_bits_cache = xbar_in_0_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_bits_cache = xbar_in_0_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_2_bits_cache = xbar_in_0_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_3_bits_cache = xbar_in_0_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_0_bits_prot = xbar_in_0_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_bits_prot = xbar_in_0_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_2_bits_prot = xbar_in_0_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_3_bits_prot = xbar_in_0_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_0_bits_qos = xbar_in_0_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_bits_qos = xbar_in_0_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_2_bits_qos = xbar_in_0_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_3_bits_qos = xbar_in_0_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_0_bits_data = xbar_in_0_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_1_bits_data = xbar_in_0_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_2_bits_data = xbar_in_0_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_3_bits_data = xbar_in_0_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_0_bits_strb = xbar_in_0_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_1_bits_strb = xbar_in_0_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_2_bits_strb = xbar_in_0_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_3_bits_strb = xbar_in_0_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_0_bits_last = xbar_in_0_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_1_bits_last = xbar_in_0_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_2_bits_last = xbar_in_0_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_3_bits_last = xbar_in_0_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  assign xbar_anonIn_b_valid = xbar_in_0_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_b_bits_resp = xbar_in_0_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_portsAROI_filtered_0_bits_id = xbar_in_0_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_bits_id = xbar_in_0_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_2_bits_id = xbar_in_0_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_3_bits_id = xbar_in_0_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_0_bits_addr = xbar_in_0_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_1_bits_addr = xbar_in_0_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_2_bits_addr = xbar_in_0_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_3_bits_addr = xbar_in_0_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_0_bits_len = xbar_in_0_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_1_bits_len = xbar_in_0_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_2_bits_len = xbar_in_0_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_3_bits_len = xbar_in_0_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_0_bits_size = xbar_in_0_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_bits_size = xbar_in_0_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_2_bits_size = xbar_in_0_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_3_bits_size = xbar_in_0_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_0_bits_burst = xbar_in_0_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_1_bits_burst = xbar_in_0_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_2_bits_burst = xbar_in_0_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_3_bits_burst = xbar_in_0_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_0_bits_lock = xbar_in_0_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_1_bits_lock = xbar_in_0_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_2_bits_lock = xbar_in_0_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_3_bits_lock = xbar_in_0_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_0_bits_cache = xbar_in_0_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_bits_cache = xbar_in_0_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_2_bits_cache = xbar_in_0_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_3_bits_cache = xbar_in_0_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_0_bits_prot = xbar_in_0_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_bits_prot = xbar_in_0_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_2_bits_prot = xbar_in_0_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_3_bits_prot = xbar_in_0_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_0_bits_qos = xbar_in_0_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_bits_qos = xbar_in_0_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_2_bits_qos = xbar_in_0_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_3_bits_qos = xbar_in_0_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  assign xbar_anonIn_r_valid = xbar_in_0_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_r_bits_data = xbar_in_0_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_r_bits_resp = xbar_in_0_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_r_bits_last = xbar_in_0_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_portsAWOI_filtered_1_0_bits_id = xbar_in_1_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_1_bits_id = xbar_in_1_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_2_bits_id = xbar_in_1_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_3_bits_id = xbar_in_1_aw_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_1_0_bits_addr = xbar_in_1_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_1_1_bits_addr = xbar_in_1_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_1_2_bits_addr = xbar_in_1_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAWOI_filtered_1_3_bits_addr = xbar_in_1_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_1_0_bits_len = xbar_in_1_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_1_1_bits_len = xbar_in_1_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_1_2_bits_len = xbar_in_1_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAWOI_filtered_1_3_bits_len = xbar_in_1_aw_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_0_bits_size = xbar_in_1_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_1_bits_size = xbar_in_1_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_2_bits_size = xbar_in_1_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_3_bits_size = xbar_in_1_aw_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_1_0_bits_burst = xbar_in_1_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_1_1_bits_burst = xbar_in_1_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_1_2_bits_burst = xbar_in_1_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAWOI_filtered_1_3_bits_burst = xbar_in_1_aw_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_1_0_bits_lock = xbar_in_1_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_1_1_bits_lock = xbar_in_1_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_1_2_bits_lock = xbar_in_1_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAWOI_filtered_1_3_bits_lock = xbar_in_1_aw_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_0_bits_cache = xbar_in_1_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_1_bits_cache = xbar_in_1_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_2_bits_cache = xbar_in_1_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_3_bits_cache = xbar_in_1_aw_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_0_bits_prot = xbar_in_1_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_1_bits_prot = xbar_in_1_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_2_bits_prot = xbar_in_1_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAWOI_filtered_1_3_bits_prot = xbar_in_1_aw_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_0_bits_qos = xbar_in_1_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_1_bits_qos = xbar_in_1_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_2_bits_qos = xbar_in_1_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAWOI_filtered_1_3_bits_qos = xbar_in_1_aw_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_1_0_bits_data = xbar_in_1_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_1_1_bits_data = xbar_in_1_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_1_2_bits_data = xbar_in_1_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [127:0] xbar_portsWOI_filtered_1_3_bits_data = xbar_in_1_w_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_1_0_bits_strb = xbar_in_1_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_1_1_bits_strb = xbar_in_1_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_1_2_bits_strb = xbar_in_1_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [15:0]  xbar_portsWOI_filtered_1_3_bits_strb = xbar_in_1_w_bits_strb;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_1_0_bits_last = xbar_in_1_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_1_1_bits_last = xbar_in_1_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_1_2_bits_last = xbar_in_1_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsWOI_filtered_1_3_bits_last = xbar_in_1_w_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  assign xbar_anonIn_1_b_valid = xbar_in_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_1_b_bits_resp = xbar_in_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  wire [2:0]   xbar_portsAROI_filtered_1_0_bits_id = xbar_in_1_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_1_bits_id = xbar_in_1_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_2_bits_id = xbar_in_1_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_3_bits_id = xbar_in_1_ar_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_1_0_bits_addr = xbar_in_1_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_1_1_bits_addr = xbar_in_1_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_1_2_bits_addr = xbar_in_1_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [29:0]  xbar_portsAROI_filtered_1_3_bits_addr = xbar_in_1_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_1_0_bits_len = xbar_in_1_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_1_1_bits_len = xbar_in_1_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_1_2_bits_len = xbar_in_1_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [7:0]   xbar_portsAROI_filtered_1_3_bits_len = xbar_in_1_ar_bits_len;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_0_bits_size = xbar_in_1_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_1_bits_size = xbar_in_1_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_2_bits_size = xbar_in_1_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_3_bits_size = xbar_in_1_ar_bits_size;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_1_0_bits_burst = xbar_in_1_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_1_1_bits_burst = xbar_in_1_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_1_2_bits_burst = xbar_in_1_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [1:0]   xbar_portsAROI_filtered_1_3_bits_burst = xbar_in_1_ar_bits_burst;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_1_0_bits_lock = xbar_in_1_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_1_1_bits_lock = xbar_in_1_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_1_2_bits_lock = xbar_in_1_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire         xbar_portsAROI_filtered_1_3_bits_lock = xbar_in_1_ar_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_0_bits_cache = xbar_in_1_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_1_bits_cache = xbar_in_1_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_2_bits_cache = xbar_in_1_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_3_bits_cache = xbar_in_1_ar_bits_cache;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_0_bits_prot = xbar_in_1_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_1_bits_prot = xbar_in_1_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_2_bits_prot = xbar_in_1_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [2:0]   xbar_portsAROI_filtered_1_3_bits_prot = xbar_in_1_ar_bits_prot;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_0_bits_qos = xbar_in_1_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_1_bits_qos = xbar_in_1_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_2_bits_qos = xbar_in_1_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  wire [3:0]   xbar_portsAROI_filtered_1_3_bits_qos = xbar_in_1_ar_bits_qos;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24
  assign xbar_anonIn_1_r_valid = xbar_in_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_1_r_bits_data = xbar_in_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_1_r_bits_resp = xbar_in_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_1_r_bits_last = xbar_in_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_in_0_aw_bits_id = {2'h2, xbar_anonIn_aw_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :103:47
  assign xbar_in_0_ar_bits_id = {2'h2, xbar_anonIn_ar_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :104:47
  wire [1:0]   xbar_arTag_lo = {xbar_requestARIO_0_1, xbar_requestARIO_0_0};	// src/main/scala/amba/axi4/Xbar.scala:77:48, :117:45
  wire [1:0]   xbar_arTag_lo_1 = xbar_arTag_lo;	// src/main/scala/amba/axi4/Xbar.scala:117:45, src/main/scala/chisel3/util/OneHot.scala:31:18
  wire [1:0]   xbar_arTag_hi = {xbar_requestARIO_0_3, xbar_requestARIO_0_2};	// src/main/scala/amba/axi4/Xbar.scala:77:48, :117:45
  wire [1:0]   xbar_arTag_hi_1 = xbar_arTag_hi;	// src/main/scala/amba/axi4/Xbar.scala:117:45, src/main/scala/chisel3/util/OneHot.scala:30:18
  wire [1:0]   xbar_arTag = {|xbar_arTag_hi_1, xbar_arTag_hi_1[1] | xbar_arTag_lo_1[1]};	// src/main/scala/chisel3/util/OneHot.scala:30:18, :31:18, :32:{10,14,28}
  wire [1:0]   xbar_awTag_lo_1 = xbar_awTag_lo;	// src/main/scala/amba/axi4/Xbar.scala:118:45, src/main/scala/chisel3/util/OneHot.scala:31:18
  wire [1:0]   xbar_awTag_hi_1 = xbar_awTag_hi;	// src/main/scala/amba/axi4/Xbar.scala:118:45, src/main/scala/chisel3/util/OneHot.scala:30:18
  wire [1:0]   xbar_awTag = {|xbar_awTag_hi_1, xbar_awTag_hi_1[1] | xbar_awTag_lo_1[1]};	// src/main/scala/chisel3/util/OneHot.scala:30:18, :31:18, :32:{10,14,28}
  wire         xbar__arFIFOMap_0_T = xbar_anonIn_ar_ready & xbar_anonIn_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/chisel3/util/Decoupled.scala:52:35
  wire         xbar__arFIFOMap_0_T_4 =
    xbar_anonIn_r_ready & xbar_anonIn_r_valid & xbar_anonIn_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:144:43, src/main/scala/chisel3/util/Decoupled.scala:52:35
  reg  [2:0]   xbar_arFIFOMap_0_count;	// src/main/scala/amba/axi4/Xbar.scala:128:34
  reg  [1:0]   xbar_arFIFOMap_0_last;	// src/main/scala/amba/axi4/Xbar.scala:129:29
  wire         xbar__arFIFOMap_0_T_12 = xbar_arFIFOMap_0_count != 3'h7;	// src/main/scala/amba/axi4/Xbar.scala:128:34, :132:43
  wire         xbar_arFIFOMap_0_portMatch = xbar_arFIFOMap_0_last == xbar_arTag;	// src/main/scala/amba/axi4/Xbar.scala:129:29, :135:71, src/main/scala/chisel3/util/OneHot.scala:32:10
  wire         xbar_arFIFOMap_0 =
    (xbar_arFIFOMap_0_count == 3'h0 | xbar_arFIFOMap_0_portMatch)
    & xbar__arFIFOMap_0_T_12;	// src/main/scala/amba/axi4/Xbar.scala:111:36, :128:34, :132:43, :135:71, :136:{22,30,44}
  wire         xbar__awFIFOMap_0_T = xbar_anonIn_aw_ready & xbar_anonIn_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/chisel3/util/Decoupled.scala:52:35
  wire         xbar__awFIFOMap_0_T_2 = xbar_anonIn_b_ready & xbar_anonIn_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/chisel3/util/Decoupled.scala:52:35
  reg  [2:0]   xbar_awFIFOMap_0_count;	// src/main/scala/amba/axi4/Xbar.scala:128:34
  reg  [1:0]   xbar_awFIFOMap_0_last;	// src/main/scala/amba/axi4/Xbar.scala:129:29
  wire         xbar__awFIFOMap_0_T_11 = xbar_awFIFOMap_0_count != 3'h7;	// src/main/scala/amba/axi4/Xbar.scala:128:34, :132:43
  wire         xbar_awFIFOMap_0_portMatch = xbar_awFIFOMap_0_last == xbar_awTag;	// src/main/scala/amba/axi4/Xbar.scala:129:29, :135:71, src/main/scala/chisel3/util/OneHot.scala:32:10
  wire         xbar_awFIFOMap_0 =
    (xbar_awFIFOMap_0_count == 3'h0 | xbar_awFIFOMap_0_portMatch)
    & xbar__awFIFOMap_0_T_11;	// src/main/scala/amba/axi4/Xbar.scala:112:36, :128:34, :132:43, :135:71, :136:{22,30,44}
  wire         xbar_in_0_ar_ready;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_ar_valid = xbar_anonIn_ar_valid & xbar_arFIFOMap_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :111:36, :153:45
  assign xbar_anonIn_ar_ready = xbar_in_0_ar_ready & xbar_arFIFOMap_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :111:36, :154:45
  reg          xbar_latched;	// src/main/scala/amba/axi4/Xbar.scala:161:30
  wire         xbar__anonIn_aw_ready_T = xbar_latched | xbar_awIn_0_io_enq_ready;	// src/main/scala/amba/axi4/Xbar.scala:161:30, :162:57
  wire         xbar_in_0_aw_ready;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_aw_valid =
    xbar_anonIn_aw_valid & xbar__anonIn_aw_ready_T & xbar_awFIFOMap_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :112:36, :162:{45,57,82}
  assign xbar_anonIn_aw_ready =
    xbar_in_0_aw_ready & xbar__anonIn_aw_ready_T & xbar_awFIFOMap_0;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :112:36, :162:57, :163:{45,82}
  assign xbar_awIn_0_io_enq_valid = xbar_anonIn_aw_valid & ~xbar_latched;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:161:30, :164:{51,54}
  wire         xbar_in_0_w_ready;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_0_w_valid = xbar_anonIn_w_valid & xbar_awIn_0_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :169:43
  assign xbar_anonIn_w_ready = xbar_in_0_w_ready & xbar_awIn_0_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :170:43
  assign xbar_awIn_0_io_deq_ready =
    xbar_anonIn_w_valid & xbar_anonIn_w_bits_last & xbar_in_0_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :171:{50,74}
  assign xbar_in_1_aw_bits_id = {1'h0, xbar_anonIn_1_aw_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :103:24
  assign xbar_in_1_ar_bits_id = {1'h0, xbar_anonIn_1_ar_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :104:24
  wire [2:0]   xbar_in_1_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_1_r_bits_id = xbar_in_1_r_bits_id[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :100:65
  wire [2:0]   xbar_in_1_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  assign xbar_anonIn_1_b_bits_id = xbar_in_1_b_bits_id[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :100:65
  wire [3:0]   xbar__arSel_T = 4'h1 << xbar_arSel_shiftAmount;	// src/main/scala/chisel3/util/OneHot.scala:64:49, :65:12
  wire [2:0]   xbar_arSel = xbar__arSel_T[2:0];	// src/main/scala/chisel3/util/OneHot.scala:65:{12,27}
  wire [3:0]   xbar__awSel_T = 4'h1 << xbar_awSel_shiftAmount;	// src/main/scala/chisel3/util/OneHot.scala:64:49, :65:12
  wire [2:0]   xbar_awSel = xbar__awSel_T[2:0];	// src/main/scala/chisel3/util/OneHot.scala:65:{12,27}
  wire [3:0]   xbar__rSel_T = 4'h1 << xbar_rSel_shiftAmount;	// src/main/scala/chisel3/util/OneHot.scala:64:49, :65:12
  wire [2:0]   xbar_rSel = xbar__rSel_T[2:0];	// src/main/scala/chisel3/util/OneHot.scala:65:{12,27}
  wire [3:0]   xbar__bSel_T = 4'h1 << xbar_bSel_shiftAmount;	// src/main/scala/chisel3/util/OneHot.scala:64:49, :65:12
  wire [2:0]   xbar_bSel = xbar__bSel_T[2:0];	// src/main/scala/chisel3/util/OneHot.scala:65:{12,27}
  wire [1:0]   xbar_arTag_lo_2 = {xbar_requestARIO_1_1, xbar_requestARIO_1_0};	// src/main/scala/amba/axi4/Xbar.scala:77:48, :117:45
  wire [1:0]   xbar_arTag_lo_3 = xbar_arTag_lo_2;	// src/main/scala/amba/axi4/Xbar.scala:117:45, src/main/scala/chisel3/util/OneHot.scala:31:18
  wire [1:0]   xbar_arTag_hi_2 = {xbar_requestARIO_1_3, xbar_requestARIO_1_2};	// src/main/scala/amba/axi4/Xbar.scala:77:48, :117:45
  wire [1:0]   xbar_arTag_hi_3 = xbar_arTag_hi_2;	// src/main/scala/amba/axi4/Xbar.scala:117:45, src/main/scala/chisel3/util/OneHot.scala:30:18
  wire [1:0]   xbar_arTag_1 = {|xbar_arTag_hi_3, xbar_arTag_hi_3[1] | xbar_arTag_lo_3[1]};	// src/main/scala/chisel3/util/OneHot.scala:30:18, :31:18, :32:{10,14,28}
  wire [1:0]   xbar_awTag_lo_3 = xbar_awTag_lo_2;	// src/main/scala/amba/axi4/Xbar.scala:118:45, src/main/scala/chisel3/util/OneHot.scala:31:18
  wire [1:0]   xbar_awTag_hi_3 = xbar_awTag_hi_2;	// src/main/scala/amba/axi4/Xbar.scala:118:45, src/main/scala/chisel3/util/OneHot.scala:30:18
  wire [1:0]   xbar_awTag_1 = {|xbar_awTag_hi_3, xbar_awTag_hi_3[1] | xbar_awTag_lo_3[1]};	// src/main/scala/chisel3/util/OneHot.scala:30:18, :31:18, :32:{10,14,28}
  wire         xbar__arFIFOMap_2_T_2 =
    xbar_arSel[2] & xbar_anonIn_1_ar_ready & xbar_anonIn_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:143:{20,25}, src/main/scala/chisel3/util/Decoupled.scala:52:35, src/main/scala/chisel3/util/OneHot.scala:65:27
  wire         xbar__arFIFOMap_2_T_6 =
    xbar_rSel[2] & xbar_anonIn_1_r_ready & xbar_anonIn_1_r_valid
    & xbar_anonIn_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:144:{19,24,43}, src/main/scala/chisel3/util/Decoupled.scala:52:35, src/main/scala/chisel3/util/OneHot.scala:65:27
  reg  [2:0]   xbar_arFIFOMap_2_count;	// src/main/scala/amba/axi4/Xbar.scala:128:34
  reg  [1:0]   xbar_arFIFOMap_2_last;	// src/main/scala/amba/axi4/Xbar.scala:129:29
  wire         xbar__arFIFOMap_2_T_14 = xbar_arFIFOMap_2_count != 3'h7;	// src/main/scala/amba/axi4/Xbar.scala:128:34, :132:43
  wire         xbar_arFIFOMap_2_portMatch = xbar_arFIFOMap_2_last == xbar_arTag_1;	// src/main/scala/amba/axi4/Xbar.scala:129:29, :135:71, src/main/scala/chisel3/util/OneHot.scala:32:10
  wire         xbar_arFIFOMap_1_2 =
    (xbar_arFIFOMap_2_count == 3'h0 | xbar_arFIFOMap_2_portMatch)
    & xbar__arFIFOMap_2_T_14;	// src/main/scala/amba/axi4/Xbar.scala:111:36, :128:34, :132:43, :135:71, :136:{22,30,44}
  wire         xbar__awFIFOMap_2_T_2 =
    xbar_awSel[2] & xbar_anonIn_1_aw_ready & xbar_anonIn_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:147:{20,25}, src/main/scala/chisel3/util/Decoupled.scala:52:35, src/main/scala/chisel3/util/OneHot.scala:65:27
  wire         xbar__awFIFOMap_2_T_5 =
    xbar_bSel[2] & xbar_anonIn_1_b_ready & xbar_anonIn_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:148:{19,24}, src/main/scala/chisel3/util/Decoupled.scala:52:35, src/main/scala/chisel3/util/OneHot.scala:65:27
  reg  [2:0]   xbar_awFIFOMap_2_count;	// src/main/scala/amba/axi4/Xbar.scala:128:34
  reg  [1:0]   xbar_awFIFOMap_2_last;	// src/main/scala/amba/axi4/Xbar.scala:129:29
  wire         xbar__awFIFOMap_2_T_13 = xbar_awFIFOMap_2_count != 3'h7;	// src/main/scala/amba/axi4/Xbar.scala:128:34, :132:43
  wire         xbar_awFIFOMap_2_portMatch = xbar_awFIFOMap_2_last == xbar_awTag_1;	// src/main/scala/amba/axi4/Xbar.scala:129:29, :135:71, src/main/scala/chisel3/util/OneHot.scala:32:10
  wire         xbar_awFIFOMap_1_2 =
    (xbar_awFIFOMap_2_count == 3'h0 | xbar_awFIFOMap_2_portMatch)
    & xbar__awFIFOMap_2_T_13;	// src/main/scala/amba/axi4/Xbar.scala:112:36, :128:34, :132:43, :135:71, :136:{22,30,44}
  wire [3:0]   _GEN_4 = {_GEN, {{xbar_arFIFOMap_1_2}, {1'h1}, {1'h1}}};	// src/main/scala/amba/axi4/Xbar.scala:111:36, :153:45
  wire         xbar_in_1_ar_ready;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_ar_valid =
    xbar_anonIn_1_ar_valid & _GEN_4[xbar_anonIn_1_ar_bits_id];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :153:45
  assign xbar_anonIn_1_ar_ready = xbar_in_1_ar_ready & _GEN_4[xbar_anonIn_1_ar_bits_id];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :153:45, :154:45
  reg          xbar_latched_1;	// src/main/scala/amba/axi4/Xbar.scala:161:30
  wire         xbar__in_1_aw_valid_T = xbar_latched_1 | xbar_awIn_1_io_enq_ready;	// src/main/scala/amba/axi4/Xbar.scala:161:30, :162:57
  wire [3:0]   _GEN_5 = {_GEN, {{xbar_awFIFOMap_1_2}, {1'h1}, {1'h1}}};	// src/main/scala/amba/axi4/Xbar.scala:112:36, :162:82
  wire         xbar_in_1_aw_ready;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_aw_valid =
    xbar_anonIn_1_aw_valid & xbar__in_1_aw_valid_T & _GEN_5[xbar_anonIn_1_aw_bits_id];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :162:{45,57,82}
  assign xbar_anonIn_1_aw_ready =
    xbar_in_1_aw_ready & xbar__in_1_aw_valid_T & _GEN_5[xbar_anonIn_1_aw_bits_id];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :162:{57,82}, :163:{45,82}
  assign xbar_awIn_1_io_enq_valid = xbar_anonIn_1_aw_valid & ~xbar_latched_1;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:161:30, :164:{51,54}
  wire         xbar_in_1_w_ready;	// src/main/scala/amba/axi4/Xbar.scala:90:18
  wire         xbar_in_1_w_valid = xbar_anonIn_1_w_valid & xbar_awIn_1_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :169:43
  assign xbar_anonIn_1_w_ready = xbar_in_1_w_ready & xbar_awIn_1_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :170:43
  assign xbar_awIn_1_io_deq_ready =
    xbar_anonIn_1_w_valid & xbar_anonIn_1_w_bits_last & xbar_in_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/amba/axi4/Xbar.scala:90:18, :171:{50,74}
  assign xbar_anonOut_aw_bits_id = xbar_out_0_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_len = xbar_out_0_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_size = xbar_out_0_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_burst = xbar_out_0_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_lock = xbar_out_0_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_cache = xbar_out_0_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_prot = xbar_out_0_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_qos = xbar_out_0_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_w_bits_data = xbar_out_0_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_w_bits_strb = xbar_out_0_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_w_bits_last = xbar_out_0_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_b_ready = xbar_out_0_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsBIO_filtered_0_bits_id = xbar_out_0_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsBIO_filtered_1_bits_id = xbar_out_0_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_0_bits_resp = xbar_out_0_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_1_bits_resp = xbar_out_0_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_anonOut_ar_valid = xbar_out_0_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_id = xbar_out_0_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_len = xbar_out_0_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_size = xbar_out_0_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_burst = xbar_out_0_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_lock = xbar_out_0_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_cache = xbar_out_0_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_prot = xbar_out_0_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_ar_bits_qos = xbar_out_0_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_r_ready = xbar_out_0_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsRIO_filtered_0_bits_id = xbar_out_0_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsRIO_filtered_1_bits_id = xbar_out_0_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_0_bits_data = xbar_out_0_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_1_bits_data = xbar_out_0_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_0_bits_resp = xbar_out_0_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_1_bits_resp = xbar_out_0_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire         xbar_portsRIO_filtered_0_bits_last = xbar_out_0_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire         xbar_portsRIO_filtered_1_bits_last = xbar_out_0_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_x1_anonOut_aw_bits_id = xbar_out_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_len = xbar_out_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_size = xbar_out_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_burst = xbar_out_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_lock = xbar_out_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_cache = xbar_out_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_prot = xbar_out_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_qos = xbar_out_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_w_bits_data = xbar_out_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_w_bits_strb = xbar_out_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_w_bits_last = xbar_out_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_b_ready = xbar_out_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsBIO_filtered_1_0_bits_id = xbar_out_1_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsBIO_filtered_1_1_bits_id = xbar_out_1_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_1_0_bits_resp = xbar_out_1_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_1_1_bits_resp = xbar_out_1_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_x1_anonOut_ar_valid = xbar_out_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_id = xbar_out_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_len = xbar_out_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_size = xbar_out_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_burst = xbar_out_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_lock = xbar_out_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_cache = xbar_out_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_prot = xbar_out_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_qos = xbar_out_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_r_ready = xbar_out_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsRIO_filtered_1_0_bits_id = xbar_out_1_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsRIO_filtered_1_1_bits_id = xbar_out_1_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_1_0_bits_data = xbar_out_1_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_1_1_bits_data = xbar_out_1_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_1_0_bits_resp = xbar_out_1_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_1_1_bits_resp = xbar_out_1_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire         xbar_portsRIO_filtered_1_0_bits_last = xbar_out_1_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire         xbar_portsRIO_filtered_1_1_bits_last = xbar_out_1_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_x1_anonOut_1_aw_bits_id = xbar_out_2_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_addr = xbar_out_2_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_len = xbar_out_2_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_size = xbar_out_2_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_burst = xbar_out_2_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_lock = xbar_out_2_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_cache = xbar_out_2_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_prot = xbar_out_2_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_bits_qos = xbar_out_2_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_w_bits_data = xbar_out_2_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_w_bits_strb = xbar_out_2_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_w_bits_last = xbar_out_2_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_b_ready = xbar_out_2_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsBIO_filtered_2_0_bits_id = xbar_out_2_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsBIO_filtered_2_1_bits_id = xbar_out_2_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_2_0_bits_resp = xbar_out_2_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_2_1_bits_resp = xbar_out_2_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_x1_anonOut_1_ar_valid = xbar_out_2_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_id = xbar_out_2_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_addr = xbar_out_2_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_len = xbar_out_2_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_size = xbar_out_2_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_burst = xbar_out_2_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_lock = xbar_out_2_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_cache = xbar_out_2_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_prot = xbar_out_2_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_ar_bits_qos = xbar_out_2_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_r_ready = xbar_out_2_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsRIO_filtered_2_0_bits_id = xbar_out_2_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsRIO_filtered_2_1_bits_id = xbar_out_2_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_2_0_bits_data = xbar_out_2_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_2_1_bits_data = xbar_out_2_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_2_0_bits_resp = xbar_out_2_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_2_1_bits_resp = xbar_out_2_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire         xbar_portsRIO_filtered_2_0_bits_last = xbar_out_2_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire         xbar_portsRIO_filtered_2_1_bits_last = xbar_out_2_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_x1_anonOut_2_aw_bits_id = xbar_out_3_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_addr = xbar_out_3_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_len = xbar_out_3_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_size = xbar_out_3_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_burst = xbar_out_3_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_lock = xbar_out_3_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_cache = xbar_out_3_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_prot = xbar_out_3_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_bits_qos = xbar_out_3_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_w_bits_data = xbar_out_3_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_w_bits_strb = xbar_out_3_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_w_bits_last = xbar_out_3_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_b_ready = xbar_out_3_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsBIO_filtered_3_0_bits_id = xbar_out_3_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsBIO_filtered_3_1_bits_id = xbar_out_3_b_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_3_0_bits_resp = xbar_out_3_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsBIO_filtered_3_1_bits_resp = xbar_out_3_b_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_x1_anonOut_2_ar_valid = xbar_out_3_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_id = xbar_out_3_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_addr = xbar_out_3_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_len = xbar_out_3_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_size = xbar_out_3_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_burst = xbar_out_3_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_lock = xbar_out_3_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_cache = xbar_out_3_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_prot = xbar_out_3_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_ar_bits_qos = xbar_out_3_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_r_ready = xbar_out_3_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19
  wire [2:0]   xbar_portsRIO_filtered_3_0_bits_id = xbar_out_3_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [2:0]   xbar_portsRIO_filtered_3_1_bits_id = xbar_out_3_r_bits_id;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_3_0_bits_data = xbar_out_3_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [127:0] xbar_portsRIO_filtered_3_1_bits_data = xbar_out_3_r_bits_data;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_3_0_bits_resp = xbar_out_3_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [1:0]   xbar_portsRIO_filtered_3_1_bits_resp = xbar_out_3_r_bits_resp;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire [29:0]  xbar_out_0_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  wire         xbar_portsRIO_filtered_3_0_bits_last = xbar_out_3_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  wire         xbar_portsRIO_filtered_3_1_bits_last = xbar_out_3_r_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24
  assign xbar_anonOut_ar_bits_addr = xbar_out_0_ar_bits_addr[27:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :182:37
  wire [29:0]  xbar_out_0_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_bits_addr = xbar_out_0_aw_bits_addr[27:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :182:37
  reg          xbar_latched_2;	// src/main/scala/amba/axi4/Xbar.scala:186:30
  wire         xbar__anonOut_aw_valid_T = xbar_latched_2 | xbar_awOut_0_io_enq_ready;	// src/main/scala/amba/axi4/Xbar.scala:186:30, :187:59
  wire         xbar_out_0_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_aw_valid = xbar_out_0_aw_valid & xbar__anonOut_aw_valid_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:{47,59}
  wire         xbar_out_0_aw_ready = xbar_anonOut_aw_ready & xbar__anonOut_aw_valid_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:59, :188:47
  assign xbar_awOut_0_io_enq_valid = xbar_out_0_aw_valid & ~xbar_latched_2;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :186:30, :189:{50,53}
  wire         xbar_out_0_w_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_anonOut_w_valid = xbar_out_0_w_valid & xbar_awOut_0_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :194:45
  wire         xbar_out_0_w_ready = xbar_anonOut_w_ready & xbar_awOut_0_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :195:45
  assign xbar_awOut_0_io_deq_ready =
    xbar_out_0_w_valid & xbar_out_0_w_bits_last & xbar_anonOut_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :196:{49,71}
  wire [29:0]  xbar_out_1_ar_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_ar_bits_addr = xbar_out_1_ar_bits_addr[28:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :182:37
  wire [29:0]  xbar_out_1_aw_bits_addr;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_bits_addr = xbar_out_1_aw_bits_addr[28:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :182:37
  reg          xbar_latched_3;	// src/main/scala/amba/axi4/Xbar.scala:186:30
  wire         xbar__out_1_aw_ready_T = xbar_latched_3 | xbar_awOut_1_io_enq_ready;	// src/main/scala/amba/axi4/Xbar.scala:186:30, :187:59
  wire         xbar_out_1_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_aw_valid = xbar_out_1_aw_valid & xbar__out_1_aw_ready_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:{47,59}
  wire         xbar_out_1_aw_ready = xbar_x1_anonOut_aw_ready & xbar__out_1_aw_ready_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:59, :188:47
  assign xbar_awOut_1_io_enq_valid = xbar_out_1_aw_valid & ~xbar_latched_3;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :186:30, :189:{50,53}
  wire         xbar_out_1_w_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_w_valid = xbar_out_1_w_valid & xbar_awOut_1_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :194:45
  wire         xbar_out_1_w_ready = xbar_x1_anonOut_w_ready & xbar_awOut_1_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :195:45
  assign xbar_awOut_1_io_deq_ready =
    xbar_out_1_w_valid & xbar_out_1_w_bits_last & xbar_x1_anonOut_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :196:{49,71}
  reg          xbar_latched_4;	// src/main/scala/amba/axi4/Xbar.scala:186:30
  wire         xbar__out_2_aw_ready_T = xbar_latched_4 | xbar_awOut_2_io_enq_ready;	// src/main/scala/amba/axi4/Xbar.scala:186:30, :187:59
  wire         xbar_out_2_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_aw_valid = xbar_out_2_aw_valid & xbar__out_2_aw_ready_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:{47,59}
  wire         xbar_out_2_aw_ready = xbar_x1_anonOut_1_aw_ready & xbar__out_2_aw_ready_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:59, :188:47
  assign xbar_awOut_2_io_enq_valid = xbar_out_2_aw_valid & ~xbar_latched_4;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :186:30, :189:{50,53}
  wire         xbar_out_2_w_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_1_w_valid = xbar_out_2_w_valid & xbar_awOut_2_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :194:45
  wire         xbar_out_2_w_ready = xbar_x1_anonOut_1_w_ready & xbar_awOut_2_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :195:45
  assign xbar_awOut_2_io_deq_ready =
    xbar_out_2_w_valid & xbar_out_2_w_bits_last & xbar_x1_anonOut_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :196:{49,71}
  reg          xbar_latched_5;	// src/main/scala/amba/axi4/Xbar.scala:186:30
  wire         xbar__out_3_aw_ready_T = xbar_latched_5 | xbar_awOut_3_io_enq_ready;	// src/main/scala/amba/axi4/Xbar.scala:186:30, :187:59
  wire         xbar_out_3_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_aw_valid = xbar_out_3_aw_valid & xbar__out_3_aw_ready_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:{47,59}
  wire         xbar_out_3_aw_ready = xbar_x1_anonOut_2_aw_ready & xbar__out_3_aw_ready_T;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :187:59, :188:47
  assign xbar_awOut_3_io_enq_valid = xbar_out_3_aw_valid & ~xbar_latched_5;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :186:30, :189:{50,53}
  wire         xbar_out_3_w_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19
  assign xbar_x1_anonOut_2_w_valid = xbar_out_3_w_valid & xbar_awOut_3_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :194:45
  wire         xbar_out_3_w_ready = xbar_x1_anonOut_2_w_ready & xbar_awOut_3_io_deq_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :195:45
  assign xbar_awOut_3_io_deq_ready =
    xbar_out_3_w_valid & xbar_out_3_w_bits_last & xbar_x1_anonOut_2_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/amba/axi4/Xbar.scala:178:19, :196:{49,71}
  wire         xbar_portsAROI_filtered_0_valid =
    xbar_in_0_ar_valid & xbar_requestARIO_0_0;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_1_valid =
    xbar_in_0_ar_valid & xbar_requestARIO_0_1;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_2_valid =
    xbar_in_0_ar_valid & xbar_requestARIO_0_2;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAROI_filtered_3_valid =
    xbar_in_0_ar_valid & xbar_requestARIO_0_3;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAROI_filtered_2_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAROI_filtered_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_in_0_ar_ready =
    xbar_requestARIO_0_0 & xbar_portsAROI_filtered_0_ready | xbar_requestARIO_0_1
    & xbar_portsAROI_filtered_1_ready | xbar_requestARIO_0_2
    & xbar_portsAROI_filtered_2_ready | xbar_requestARIO_0_3
    & xbar_portsAROI_filtered_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73
  wire         xbar_portsAROI_filtered_1_0_valid =
    xbar_in_1_ar_valid & xbar_requestARIO_1_0;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_1_1_valid =
    xbar_in_1_ar_valid & xbar_requestARIO_1_1;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_1_2_valid =
    xbar_in_1_ar_valid & xbar_requestARIO_1_2;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_1_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAROI_filtered_1_3_valid =
    xbar_in_1_ar_valid & xbar_requestARIO_1_3;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, :252:40
  wire         xbar_portsAROI_filtered_1_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAROI_filtered_1_2_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAROI_filtered_1_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_in_1_ar_ready =
    xbar_requestARIO_1_0 & xbar_portsAROI_filtered_1_0_ready | xbar_requestARIO_1_1
    & xbar_portsAROI_filtered_1_1_ready | xbar_requestARIO_1_2
    & xbar_portsAROI_filtered_1_2_ready | xbar_requestARIO_1_3
    & xbar_portsAROI_filtered_1_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:77:48, :90:18, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73
  wire         xbar_portsAWOI_filtered_0_valid =
    xbar_in_0_aw_valid & xbar_requestAWIO_0_0;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_1_valid =
    xbar_in_0_aw_valid & xbar_requestAWIO_0_1;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_2_valid =
    xbar_in_0_aw_valid & xbar_requestAWIO_0_2;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAWOI_filtered_3_valid =
    xbar_in_0_aw_valid & xbar_requestAWIO_0_3;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAWOI_filtered_2_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAWOI_filtered_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_in_0_aw_ready =
    xbar_requestAWIO_0_0 & xbar_portsAWOI_filtered_0_ready | xbar_requestAWIO_0_1
    & xbar_portsAWOI_filtered_1_ready | xbar_requestAWIO_0_2
    & xbar_portsAWOI_filtered_2_ready | xbar_requestAWIO_0_3
    & xbar_portsAWOI_filtered_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73
  wire         xbar_portsAWOI_filtered_1_0_valid =
    xbar_in_1_aw_valid & xbar_requestAWIO_1_0;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_1_1_valid =
    xbar_in_1_aw_valid & xbar_requestAWIO_1_1;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_1_2_valid =
    xbar_in_1_aw_valid & xbar_requestAWIO_1_2;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_1_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAWOI_filtered_1_3_valid =
    xbar_in_1_aw_valid & xbar_requestAWIO_1_3;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, :252:40
  wire         xbar_portsAWOI_filtered_1_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAWOI_filtered_1_2_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsAWOI_filtered_1_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_in_1_aw_ready =
    xbar_requestAWIO_1_0 & xbar_portsAWOI_filtered_1_0_ready | xbar_requestAWIO_1_1
    & xbar_portsAWOI_filtered_1_1_ready | xbar_requestAWIO_1_2
    & xbar_portsAWOI_filtered_1_2_ready | xbar_requestAWIO_1_3
    & xbar_portsAWOI_filtered_1_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:78:48, :90:18, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73
  wire         xbar_portsWOI_filtered_0_valid = xbar_in_0_w_valid & xbar_requestWIO_0_0;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_1_valid = xbar_in_0_w_valid & xbar_requestWIO_0_1;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_2_valid = xbar_in_0_w_valid & xbar_requestWIO_0_2;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsWOI_filtered_3_valid = xbar_in_0_w_valid & xbar_requestWIO_0_3;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsWOI_filtered_2_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsWOI_filtered_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_in_0_w_ready =
    xbar_requestWIO_0_0 & xbar_portsWOI_filtered_0_ready | xbar_requestWIO_0_1
    & xbar_portsWOI_filtered_1_ready | xbar_requestWIO_0_2
    & xbar_portsWOI_filtered_2_ready | xbar_requestWIO_0_3
    & xbar_portsWOI_filtered_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73
  wire         xbar_portsWOI_filtered_1_0_valid = xbar_in_1_w_valid & xbar_requestWIO_1_0;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_1_1_valid = xbar_in_1_w_valid & xbar_requestWIO_1_1;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_1_2_valid = xbar_in_1_w_valid & xbar_requestWIO_1_2;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_1_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsWOI_filtered_1_3_valid = xbar_in_1_w_valid & xbar_requestWIO_1_3;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, :252:40
  wire         xbar_portsWOI_filtered_1_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsWOI_filtered_1_2_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsWOI_filtered_1_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_in_1_w_ready =
    xbar_requestWIO_1_0 & xbar_portsWOI_filtered_1_0_ready | xbar_requestWIO_1_1
    & xbar_portsWOI_filtered_1_1_ready | xbar_requestWIO_1_2
    & xbar_portsWOI_filtered_1_2_ready | xbar_requestWIO_1_3
    & xbar_portsWOI_filtered_1_3_ready;	// src/main/scala/amba/axi4/Xbar.scala:84:73, :90:18, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73
  wire         xbar_portsRIO_filtered_0_valid = xbar_out_0_r_valid & xbar_requestROI_0_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsRIO_filtered_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsRIO_filtered_1_valid = xbar_out_0_r_valid & xbar_requestROI_0_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsRIO_filtered_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_0_r_ready =
    xbar_requestROI_0_0 & xbar_portsRIO_filtered_0_ready | xbar_requestROI_0_1
    & xbar_portsRIO_filtered_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  wire         xbar_portsRIO_filtered_1_0_valid =
    xbar_out_1_r_valid & xbar_requestROI_1_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsRIO_filtered_1_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsRIO_filtered_1_1_valid =
    xbar_out_1_r_valid & xbar_requestROI_1_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsRIO_filtered_1_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_1_r_ready =
    xbar_requestROI_1_0 & xbar_portsRIO_filtered_1_0_ready | xbar_requestROI_1_1
    & xbar_portsRIO_filtered_1_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  wire         xbar_portsRIO_filtered_2_0_valid =
    xbar_out_2_r_valid & xbar_requestROI_2_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsRIO_filtered_2_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsRIO_filtered_2_1_valid =
    xbar_out_2_r_valid & xbar_requestROI_2_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsRIO_filtered_2_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_2_r_ready =
    xbar_requestROI_2_0 & xbar_portsRIO_filtered_2_0_ready | xbar_requestROI_2_1
    & xbar_portsRIO_filtered_2_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  wire         xbar_portsRIO_filtered_3_0_valid =
    xbar_out_3_r_valid & xbar_requestROI_3_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsRIO_filtered_3_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsRIO_filtered_3_1_valid =
    xbar_out_3_r_valid & xbar_requestROI_3_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsRIO_filtered_3_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_3_r_ready =
    xbar_requestROI_3_0 & xbar_portsRIO_filtered_3_0_ready | xbar_requestROI_3_1
    & xbar_portsRIO_filtered_3_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  wire         xbar_portsBIO_filtered_0_valid = xbar_out_0_b_valid & xbar_requestBOI_0_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsBIO_filtered_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsBIO_filtered_1_valid = xbar_out_0_b_valid & xbar_requestBOI_0_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsBIO_filtered_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_0_b_ready =
    xbar_requestBOI_0_0 & xbar_portsBIO_filtered_0_ready | xbar_requestBOI_0_1
    & xbar_portsBIO_filtered_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  wire         xbar_portsBIO_filtered_1_0_valid =
    xbar_out_1_b_valid & xbar_requestBOI_1_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsBIO_filtered_1_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsBIO_filtered_1_1_valid =
    xbar_out_1_b_valid & xbar_requestBOI_1_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsBIO_filtered_1_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_1_b_ready =
    xbar_requestBOI_1_0 & xbar_portsBIO_filtered_1_0_ready | xbar_requestBOI_1_1
    & xbar_portsBIO_filtered_1_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  wire         xbar_portsBIO_filtered_2_0_valid =
    xbar_out_2_b_valid & xbar_requestBOI_2_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsBIO_filtered_2_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsBIO_filtered_2_1_valid =
    xbar_out_2_b_valid & xbar_requestBOI_2_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsBIO_filtered_2_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_2_b_ready =
    xbar_requestBOI_2_0 & xbar_portsBIO_filtered_2_0_ready | xbar_requestBOI_2_1
    & xbar_portsBIO_filtered_2_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  wire         xbar_portsBIO_filtered_3_0_valid =
    xbar_out_3_b_valid & xbar_requestBOI_3_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:46:9
  wire         xbar_portsBIO_filtered_3_0_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  wire         xbar_portsBIO_filtered_3_1_valid =
    xbar_out_3_b_valid & xbar_requestBOI_3_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :252:40, src/main/scala/diplomacy/Parameters.scala:56:48
  wire         xbar_portsBIO_filtered_3_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:249:24
  assign xbar_out_3_b_ready =
    xbar_requestBOI_3_0 & xbar_portsBIO_filtered_3_0_ready | xbar_requestBOI_3_1
    & xbar_portsBIO_filtered_3_1_ready;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, src/main/scala/diplomacy/Parameters.scala:46:9, :56:48
  reg          xbar_awOut_0_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_awOut_0_io_enq_bits_anyValid =
    xbar_portsAWOI_filtered_0_valid | xbar_portsAWOI_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_awOut_0_io_enq_bits_readys_valid =
    {xbar_portsAWOI_filtered_1_0_valid, xbar_portsAWOI_filtered_0_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_awOut_0_io_enq_bits_readys_mask;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_awOut_0_io_enq_bits_readys_filter =
    {xbar_awOut_0_io_enq_bits_readys_valid & ~xbar_awOut_0_io_enq_bits_readys_mask,
     xbar_awOut_0_io_enq_bits_readys_valid};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_awOut_0_io_enq_bits_readys_unready =
    {xbar_awOut_0_io_enq_bits_readys_mask[1],
     xbar_awOut_0_io_enq_bits_readys_filter[3] | xbar_awOut_0_io_enq_bits_readys_mask[0],
     xbar_awOut_0_io_enq_bits_readys_filter[2:1]
       | xbar_awOut_0_io_enq_bits_readys_filter[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_awOut_0_io_enq_bits_readys_readys =
    ~(xbar_awOut_0_io_enq_bits_readys_unready[3:2]
      & xbar_awOut_0_io_enq_bits_readys_unready[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_awOut_0_io_enq_bits_readys_0 =
    xbar_awOut_0_io_enq_bits_readys_readys[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_0_io_enq_bits_readys_1 =
    xbar_awOut_0_io_enq_bits_readys_readys[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_0_io_enq_bits_winner_0 =
    xbar_awOut_0_io_enq_bits_readys_0 & xbar_portsAWOI_filtered_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_0_io_enq_bits_winner_1 =
    xbar_awOut_0_io_enq_bits_readys_1 & xbar_portsAWOI_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_0_io_enq_bits_prefixOR_1 = xbar_awOut_0_io_enq_bits_winner_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_awOut_0_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_awOut_0_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_awOut_0_io_enq_bits_muxState_0 =
    xbar_awOut_0_io_enq_bits_idle
      ? xbar_awOut_0_io_enq_bits_winner_0
      : xbar_awOut_0_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_0_io_enq_bits_muxState_1 =
    xbar_awOut_0_io_enq_bits_idle
      ? xbar_awOut_0_io_enq_bits_winner_1
      : xbar_awOut_0_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_0_io_enq_bits_allowed_0 =
    xbar_awOut_0_io_enq_bits_idle
      ? xbar_awOut_0_io_enq_bits_readys_0
      : xbar_awOut_0_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_awOut_0_io_enq_bits_allowed_1 =
    xbar_awOut_0_io_enq_bits_idle
      ? xbar_awOut_0_io_enq_bits_readys_1
      : xbar_awOut_0_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAWOI_filtered_0_ready =
    xbar_out_0_aw_ready & xbar_awOut_0_io_enq_bits_allowed_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAWOI_filtered_1_0_ready =
    xbar_out_0_aw_ready & xbar_awOut_0_io_enq_bits_allowed_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_0_aw_valid =
    xbar_awOut_0_io_enq_bits_idle
      ? xbar_awOut_0_io_enq_bits_anyValid
      : xbar_awOut_0_io_enq_bits_state_0 & xbar_portsAWOI_filtered_0_valid
        | xbar_awOut_0_io_enq_bits_state_1 & xbar_portsAWOI_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_qos =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_qos : 4'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_0_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_prot =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_prot : 3'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_0_bits_prot
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_cache =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_cache : 4'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_0_bits_cache
         : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_lock =
    xbar_awOut_0_io_enq_bits_muxState_0 & xbar_portsAWOI_filtered_0_bits_lock
    | xbar_awOut_0_io_enq_bits_muxState_1 & xbar_portsAWOI_filtered_1_0_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_burst =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_burst : 2'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_0_bits_burst
         : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_size =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_size : 3'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_0_bits_size
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_len =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_len : 8'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_0_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_addr =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_addr : 30'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_0_bits_addr
         : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_aw_bits_id =
    (xbar_awOut_0_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_0_bits_id : 3'h0)
    | (xbar_awOut_0_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_0_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_awOut_0_io_enq_bits =
    {xbar_awOut_0_io_enq_bits_muxState_1, xbar_awOut_0_io_enq_bits_muxState_0};	// src/main/scala/amba/axi4/Xbar.scala:213:81, :292:23
  reg          xbar_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid =
    xbar_portsAROI_filtered_0_valid | xbar_portsAROI_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_valid =
    {xbar_portsAROI_filtered_1_0_valid, xbar_portsAROI_filtered_0_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_readys_mask;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_readys_filter =
    {xbar_readys_valid & ~xbar_readys_mask, xbar_readys_valid};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_readys_unready =
    {xbar_readys_mask[1],
     xbar_readys_filter[3] | xbar_readys_mask[0],
     xbar_readys_filter[2:1] | xbar_readys_filter[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_readys_readys =
    ~(xbar_readys_unready[3:2] & xbar_readys_unready[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_0 = xbar_readys_readys[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_1 = xbar_readys_readys[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_0 = xbar_readys_0 & xbar_portsAROI_filtered_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_1 = xbar_readys_1 & xbar_portsAROI_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1 = xbar_winner_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_state_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_0 = xbar_idle ? xbar_winner_0 : xbar_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_1 = xbar_idle ? xbar_winner_1 : xbar_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_0 = xbar_idle ? xbar_readys_0 : xbar_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_1 = xbar_idle ? xbar_readys_1 : xbar_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAROI_filtered_0_ready = xbar_out_0_ar_ready & xbar_allowed_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAROI_filtered_1_0_ready = xbar_out_0_ar_ready & xbar_allowed_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_0_ar_valid =
    xbar_idle
      ? xbar_anyValid
      : xbar_state_0 & xbar_portsAROI_filtered_0_valid | xbar_state_1
        & xbar_portsAROI_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_qos =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_qos : 4'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_prot =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_prot : 3'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_prot : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_cache =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_cache : 4'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_cache : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_lock =
    xbar_muxState_0 & xbar_portsAROI_filtered_0_bits_lock | xbar_muxState_1
    & xbar_portsAROI_filtered_1_0_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_burst =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_burst : 2'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_burst : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_size =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_size : 3'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_size : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_len =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_len : 8'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_addr =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_addr : 30'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_addr : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_ar_bits_id =
    (xbar_muxState_0 ? xbar_portsAROI_filtered_0_bits_id : 3'h0)
    | (xbar_muxState_1 ? xbar_portsAROI_filtered_1_0_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_0_w_valid =
    xbar_awOut_0_io_deq_bits[0] & xbar_portsWOI_filtered_0_valid
    | xbar_awOut_0_io_deq_bits[1] & xbar_portsWOI_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_0_w_bits_last =
    xbar_awOut_0_io_deq_bits[0] & xbar_portsWOI_filtered_0_bits_last
    | xbar_awOut_0_io_deq_bits[1] & xbar_portsWOI_filtered_1_0_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_0_w_bits_strb =
    (xbar_awOut_0_io_deq_bits[0] ? xbar_portsWOI_filtered_0_bits_strb : 16'h0)
    | (xbar_awOut_0_io_deq_bits[1] ? xbar_portsWOI_filtered_1_0_bits_strb : 16'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_0_w_bits_data =
    (xbar_awOut_0_io_deq_bits[0] ? xbar_portsWOI_filtered_0_bits_data : 128'h0)
    | (xbar_awOut_0_io_deq_bits[1] ? xbar_portsWOI_filtered_1_0_bits_data : 128'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_portsWOI_filtered_0_ready =
    xbar_out_0_w_ready & xbar_awOut_0_io_deq_bits[0];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  assign xbar_portsWOI_filtered_1_0_ready =
    xbar_out_0_w_ready & xbar_awOut_0_io_deq_bits[1];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  reg          xbar_awOut_1_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_awOut_1_io_enq_bits_anyValid =
    xbar_portsAWOI_filtered_1_valid | xbar_portsAWOI_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_awOut_1_io_enq_bits_readys_valid =
    {xbar_portsAWOI_filtered_1_1_valid, xbar_portsAWOI_filtered_1_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_awOut_1_io_enq_bits_readys_mask;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_awOut_1_io_enq_bits_readys_filter =
    {xbar_awOut_1_io_enq_bits_readys_valid & ~xbar_awOut_1_io_enq_bits_readys_mask,
     xbar_awOut_1_io_enq_bits_readys_valid};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_awOut_1_io_enq_bits_readys_unready =
    {xbar_awOut_1_io_enq_bits_readys_mask[1],
     xbar_awOut_1_io_enq_bits_readys_filter[3] | xbar_awOut_1_io_enq_bits_readys_mask[0],
     xbar_awOut_1_io_enq_bits_readys_filter[2:1]
       | xbar_awOut_1_io_enq_bits_readys_filter[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_awOut_1_io_enq_bits_readys_readys =
    ~(xbar_awOut_1_io_enq_bits_readys_unready[3:2]
      & xbar_awOut_1_io_enq_bits_readys_unready[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_awOut_1_io_enq_bits_readys_0 =
    xbar_awOut_1_io_enq_bits_readys_readys[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_1_io_enq_bits_readys_1 =
    xbar_awOut_1_io_enq_bits_readys_readys[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_1_io_enq_bits_winner_0 =
    xbar_awOut_1_io_enq_bits_readys_0 & xbar_portsAWOI_filtered_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_1_io_enq_bits_winner_1 =
    xbar_awOut_1_io_enq_bits_readys_1 & xbar_portsAWOI_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_1_io_enq_bits_prefixOR_1 = xbar_awOut_1_io_enq_bits_winner_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_awOut_1_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_awOut_1_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_awOut_1_io_enq_bits_muxState_0 =
    xbar_awOut_1_io_enq_bits_idle
      ? xbar_awOut_1_io_enq_bits_winner_0
      : xbar_awOut_1_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_1_io_enq_bits_muxState_1 =
    xbar_awOut_1_io_enq_bits_idle
      ? xbar_awOut_1_io_enq_bits_winner_1
      : xbar_awOut_1_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_1_io_enq_bits_allowed_0 =
    xbar_awOut_1_io_enq_bits_idle
      ? xbar_awOut_1_io_enq_bits_readys_0
      : xbar_awOut_1_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_awOut_1_io_enq_bits_allowed_1 =
    xbar_awOut_1_io_enq_bits_idle
      ? xbar_awOut_1_io_enq_bits_readys_1
      : xbar_awOut_1_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAWOI_filtered_1_ready =
    xbar_out_1_aw_ready & xbar_awOut_1_io_enq_bits_allowed_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAWOI_filtered_1_1_ready =
    xbar_out_1_aw_ready & xbar_awOut_1_io_enq_bits_allowed_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_1_aw_valid =
    xbar_awOut_1_io_enq_bits_idle
      ? xbar_awOut_1_io_enq_bits_anyValid
      : xbar_awOut_1_io_enq_bits_state_0 & xbar_portsAWOI_filtered_1_valid
        | xbar_awOut_1_io_enq_bits_state_1 & xbar_portsAWOI_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_qos =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_qos : 4'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_1_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_prot =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_prot : 3'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_1_bits_prot
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_cache =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_cache : 4'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_1_bits_cache
         : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_lock =
    xbar_awOut_1_io_enq_bits_muxState_0 & xbar_portsAWOI_filtered_1_bits_lock
    | xbar_awOut_1_io_enq_bits_muxState_1 & xbar_portsAWOI_filtered_1_1_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_burst =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_burst : 2'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_1_bits_burst
         : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_size =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_size : 3'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_1_bits_size
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_len =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_len : 8'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_1_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_addr =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_addr : 30'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_1_bits_addr
         : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_aw_bits_id =
    (xbar_awOut_1_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_1_bits_id : 3'h0)
    | (xbar_awOut_1_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_1_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_awOut_1_io_enq_bits =
    {xbar_awOut_1_io_enq_bits_muxState_1, xbar_awOut_1_io_enq_bits_muxState_0};	// src/main/scala/amba/axi4/Xbar.scala:213:81, :292:23
  reg          xbar_idle_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid_1 =
    xbar_portsAROI_filtered_1_valid | xbar_portsAROI_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_valid_1 =
    {xbar_portsAROI_filtered_1_1_valid, xbar_portsAROI_filtered_1_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_readys_mask_1;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_readys_filter_1 =
    {xbar_readys_valid_1 & ~xbar_readys_mask_1, xbar_readys_valid_1};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_readys_unready_1 =
    {xbar_readys_mask_1[1],
     xbar_readys_filter_1[3] | xbar_readys_mask_1[0],
     xbar_readys_filter_1[2:1] | xbar_readys_filter_1[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_readys_readys_1 =
    ~(xbar_readys_unready_1[3:2] & xbar_readys_unready_1[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_1_0 = xbar_readys_readys_1[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_1_1 = xbar_readys_readys_1[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_1_0 = xbar_readys_1_0 & xbar_portsAROI_filtered_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_1_1 = xbar_readys_1_1 & xbar_portsAROI_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1_1 = xbar_winner_1_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_state_1_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_1_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_1_0 = xbar_idle_1 ? xbar_winner_1_0 : xbar_state_1_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_1_1 = xbar_idle_1 ? xbar_winner_1_1 : xbar_state_1_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_1_0 = xbar_idle_1 ? xbar_readys_1_0 : xbar_state_1_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_1_1 = xbar_idle_1 ? xbar_readys_1_1 : xbar_state_1_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAROI_filtered_1_ready = xbar_out_1_ar_ready & xbar_allowed_1_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAROI_filtered_1_1_ready = xbar_out_1_ar_ready & xbar_allowed_1_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_1_ar_valid =
    xbar_idle_1
      ? xbar_anyValid_1
      : xbar_state_1_0 & xbar_portsAROI_filtered_1_valid | xbar_state_1_1
        & xbar_portsAROI_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_qos =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_qos : 4'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_prot =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_prot : 3'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_prot : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_cache =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_cache : 4'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_cache : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_lock =
    xbar_muxState_1_0 & xbar_portsAROI_filtered_1_bits_lock | xbar_muxState_1_1
    & xbar_portsAROI_filtered_1_1_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_burst =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_burst : 2'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_burst : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_size =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_size : 3'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_size : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_len =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_len : 8'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_addr =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_addr : 30'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_addr : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_ar_bits_id =
    (xbar_muxState_1_0 ? xbar_portsAROI_filtered_1_bits_id : 3'h0)
    | (xbar_muxState_1_1 ? xbar_portsAROI_filtered_1_1_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_1_w_valid =
    xbar_awOut_1_io_deq_bits[0] & xbar_portsWOI_filtered_1_valid
    | xbar_awOut_1_io_deq_bits[1] & xbar_portsWOI_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_1_w_bits_last =
    xbar_awOut_1_io_deq_bits[0] & xbar_portsWOI_filtered_1_bits_last
    | xbar_awOut_1_io_deq_bits[1] & xbar_portsWOI_filtered_1_1_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_1_w_bits_strb =
    (xbar_awOut_1_io_deq_bits[0] ? xbar_portsWOI_filtered_1_bits_strb : 16'h0)
    | (xbar_awOut_1_io_deq_bits[1] ? xbar_portsWOI_filtered_1_1_bits_strb : 16'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_1_w_bits_data =
    (xbar_awOut_1_io_deq_bits[0] ? xbar_portsWOI_filtered_1_bits_data : 128'h0)
    | (xbar_awOut_1_io_deq_bits[1] ? xbar_portsWOI_filtered_1_1_bits_data : 128'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_portsWOI_filtered_1_ready =
    xbar_out_1_w_ready & xbar_awOut_1_io_deq_bits[0];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  assign xbar_portsWOI_filtered_1_1_ready =
    xbar_out_1_w_ready & xbar_awOut_1_io_deq_bits[1];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  reg          xbar_awOut_2_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_awOut_2_io_enq_bits_anyValid =
    xbar_portsAWOI_filtered_2_valid | xbar_portsAWOI_filtered_1_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_awOut_2_io_enq_bits_readys_valid =
    {xbar_portsAWOI_filtered_1_2_valid, xbar_portsAWOI_filtered_2_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_awOut_2_io_enq_bits_readys_mask;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_awOut_2_io_enq_bits_readys_filter =
    {xbar_awOut_2_io_enq_bits_readys_valid & ~xbar_awOut_2_io_enq_bits_readys_mask,
     xbar_awOut_2_io_enq_bits_readys_valid};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_awOut_2_io_enq_bits_readys_unready =
    {xbar_awOut_2_io_enq_bits_readys_mask[1],
     xbar_awOut_2_io_enq_bits_readys_filter[3] | xbar_awOut_2_io_enq_bits_readys_mask[0],
     xbar_awOut_2_io_enq_bits_readys_filter[2:1]
       | xbar_awOut_2_io_enq_bits_readys_filter[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_awOut_2_io_enq_bits_readys_readys =
    ~(xbar_awOut_2_io_enq_bits_readys_unready[3:2]
      & xbar_awOut_2_io_enq_bits_readys_unready[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_awOut_2_io_enq_bits_readys_0 =
    xbar_awOut_2_io_enq_bits_readys_readys[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_2_io_enq_bits_readys_1 =
    xbar_awOut_2_io_enq_bits_readys_readys[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_2_io_enq_bits_winner_0 =
    xbar_awOut_2_io_enq_bits_readys_0 & xbar_portsAWOI_filtered_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_2_io_enq_bits_winner_1 =
    xbar_awOut_2_io_enq_bits_readys_1 & xbar_portsAWOI_filtered_1_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_2_io_enq_bits_prefixOR_1 = xbar_awOut_2_io_enq_bits_winner_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_awOut_2_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_awOut_2_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_awOut_2_io_enq_bits_muxState_0 =
    xbar_awOut_2_io_enq_bits_idle
      ? xbar_awOut_2_io_enq_bits_winner_0
      : xbar_awOut_2_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_2_io_enq_bits_muxState_1 =
    xbar_awOut_2_io_enq_bits_idle
      ? xbar_awOut_2_io_enq_bits_winner_1
      : xbar_awOut_2_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_2_io_enq_bits_allowed_0 =
    xbar_awOut_2_io_enq_bits_idle
      ? xbar_awOut_2_io_enq_bits_readys_0
      : xbar_awOut_2_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_awOut_2_io_enq_bits_allowed_1 =
    xbar_awOut_2_io_enq_bits_idle
      ? xbar_awOut_2_io_enq_bits_readys_1
      : xbar_awOut_2_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAWOI_filtered_2_ready =
    xbar_out_2_aw_ready & xbar_awOut_2_io_enq_bits_allowed_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAWOI_filtered_1_2_ready =
    xbar_out_2_aw_ready & xbar_awOut_2_io_enq_bits_allowed_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_2_aw_valid =
    xbar_awOut_2_io_enq_bits_idle
      ? xbar_awOut_2_io_enq_bits_anyValid
      : xbar_awOut_2_io_enq_bits_state_0 & xbar_portsAWOI_filtered_2_valid
        | xbar_awOut_2_io_enq_bits_state_1 & xbar_portsAWOI_filtered_1_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_qos =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_qos : 4'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_2_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_prot =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_prot : 3'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_2_bits_prot
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_cache =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_cache : 4'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_2_bits_cache
         : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_lock =
    xbar_awOut_2_io_enq_bits_muxState_0 & xbar_portsAWOI_filtered_2_bits_lock
    | xbar_awOut_2_io_enq_bits_muxState_1 & xbar_portsAWOI_filtered_1_2_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_burst =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_burst : 2'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_2_bits_burst
         : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_size =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_size : 3'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_2_bits_size
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_len =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_len : 8'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_2_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_addr =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_addr : 30'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_2_bits_addr
         : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_aw_bits_id =
    (xbar_awOut_2_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_2_bits_id : 3'h0)
    | (xbar_awOut_2_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_2_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_awOut_2_io_enq_bits =
    {xbar_awOut_2_io_enq_bits_muxState_1, xbar_awOut_2_io_enq_bits_muxState_0};	// src/main/scala/amba/axi4/Xbar.scala:213:81, :292:23
  reg          xbar_idle_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid_2 =
    xbar_portsAROI_filtered_2_valid | xbar_portsAROI_filtered_1_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_valid_2 =
    {xbar_portsAROI_filtered_1_2_valid, xbar_portsAROI_filtered_2_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_readys_mask_2;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_readys_filter_2 =
    {xbar_readys_valid_2 & ~xbar_readys_mask_2, xbar_readys_valid_2};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_readys_unready_2 =
    {xbar_readys_mask_2[1],
     xbar_readys_filter_2[3] | xbar_readys_mask_2[0],
     xbar_readys_filter_2[2:1] | xbar_readys_filter_2[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_readys_readys_2 =
    ~(xbar_readys_unready_2[3:2] & xbar_readys_unready_2[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_2_0 = xbar_readys_readys_2[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_2_1 = xbar_readys_readys_2[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_2_0 = xbar_readys_2_0 & xbar_portsAROI_filtered_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_2_1 = xbar_readys_2_1 & xbar_portsAROI_filtered_1_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1_2 = xbar_winner_2_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_state_2_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_2_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_2_0 = xbar_idle_2 ? xbar_winner_2_0 : xbar_state_2_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_2_1 = xbar_idle_2 ? xbar_winner_2_1 : xbar_state_2_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_2_0 = xbar_idle_2 ? xbar_readys_2_0 : xbar_state_2_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_2_1 = xbar_idle_2 ? xbar_readys_2_1 : xbar_state_2_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAROI_filtered_2_ready = xbar_out_2_ar_ready & xbar_allowed_2_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAROI_filtered_1_2_ready = xbar_out_2_ar_ready & xbar_allowed_2_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_2_ar_valid =
    xbar_idle_2
      ? xbar_anyValid_2
      : xbar_state_2_0 & xbar_portsAROI_filtered_2_valid | xbar_state_2_1
        & xbar_portsAROI_filtered_1_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_qos =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_qos : 4'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_prot =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_prot : 3'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_prot : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_cache =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_cache : 4'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_cache : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_lock =
    xbar_muxState_2_0 & xbar_portsAROI_filtered_2_bits_lock | xbar_muxState_2_1
    & xbar_portsAROI_filtered_1_2_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_burst =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_burst : 2'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_burst : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_size =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_size : 3'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_size : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_len =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_len : 8'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_addr =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_addr : 30'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_addr : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_ar_bits_id =
    (xbar_muxState_2_0 ? xbar_portsAROI_filtered_2_bits_id : 3'h0)
    | (xbar_muxState_2_1 ? xbar_portsAROI_filtered_1_2_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_2_w_valid =
    xbar_awOut_2_io_deq_bits[0] & xbar_portsWOI_filtered_2_valid
    | xbar_awOut_2_io_deq_bits[1] & xbar_portsWOI_filtered_1_2_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_2_w_bits_last =
    xbar_awOut_2_io_deq_bits[0] & xbar_portsWOI_filtered_2_bits_last
    | xbar_awOut_2_io_deq_bits[1] & xbar_portsWOI_filtered_1_2_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_2_w_bits_strb =
    (xbar_awOut_2_io_deq_bits[0] ? xbar_portsWOI_filtered_2_bits_strb : 16'h0)
    | (xbar_awOut_2_io_deq_bits[1] ? xbar_portsWOI_filtered_1_2_bits_strb : 16'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_2_w_bits_data =
    (xbar_awOut_2_io_deq_bits[0] ? xbar_portsWOI_filtered_2_bits_data : 128'h0)
    | (xbar_awOut_2_io_deq_bits[1] ? xbar_portsWOI_filtered_1_2_bits_data : 128'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_portsWOI_filtered_2_ready =
    xbar_out_2_w_ready & xbar_awOut_2_io_deq_bits[0];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  assign xbar_portsWOI_filtered_1_2_ready =
    xbar_out_2_w_ready & xbar_awOut_2_io_deq_bits[1];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  reg          xbar_awOut_3_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_awOut_3_io_enq_bits_anyValid =
    xbar_portsAWOI_filtered_3_valid | xbar_portsAWOI_filtered_1_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_awOut_3_io_enq_bits_readys_valid =
    {xbar_portsAWOI_filtered_1_3_valid, xbar_portsAWOI_filtered_3_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_awOut_3_io_enq_bits_readys_mask;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_awOut_3_io_enq_bits_readys_filter =
    {xbar_awOut_3_io_enq_bits_readys_valid & ~xbar_awOut_3_io_enq_bits_readys_mask,
     xbar_awOut_3_io_enq_bits_readys_valid};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_awOut_3_io_enq_bits_readys_unready =
    {xbar_awOut_3_io_enq_bits_readys_mask[1],
     xbar_awOut_3_io_enq_bits_readys_filter[3] | xbar_awOut_3_io_enq_bits_readys_mask[0],
     xbar_awOut_3_io_enq_bits_readys_filter[2:1]
       | xbar_awOut_3_io_enq_bits_readys_filter[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_awOut_3_io_enq_bits_readys_readys =
    ~(xbar_awOut_3_io_enq_bits_readys_unready[3:2]
      & xbar_awOut_3_io_enq_bits_readys_unready[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_awOut_3_io_enq_bits_readys_0 =
    xbar_awOut_3_io_enq_bits_readys_readys[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_3_io_enq_bits_readys_1 =
    xbar_awOut_3_io_enq_bits_readys_readys[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_awOut_3_io_enq_bits_winner_0 =
    xbar_awOut_3_io_enq_bits_readys_0 & xbar_portsAWOI_filtered_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_3_io_enq_bits_winner_1 =
    xbar_awOut_3_io_enq_bits_readys_1 & xbar_portsAWOI_filtered_1_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_awOut_3_io_enq_bits_prefixOR_1 = xbar_awOut_3_io_enq_bits_winner_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_awOut_3_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_awOut_3_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_awOut_3_io_enq_bits_muxState_0 =
    xbar_awOut_3_io_enq_bits_idle
      ? xbar_awOut_3_io_enq_bits_winner_0
      : xbar_awOut_3_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_3_io_enq_bits_muxState_1 =
    xbar_awOut_3_io_enq_bits_idle
      ? xbar_awOut_3_io_enq_bits_winner_1
      : xbar_awOut_3_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_awOut_3_io_enq_bits_allowed_0 =
    xbar_awOut_3_io_enq_bits_idle
      ? xbar_awOut_3_io_enq_bits_readys_0
      : xbar_awOut_3_io_enq_bits_state_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_awOut_3_io_enq_bits_allowed_1 =
    xbar_awOut_3_io_enq_bits_idle
      ? xbar_awOut_3_io_enq_bits_readys_1
      : xbar_awOut_3_io_enq_bits_state_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAWOI_filtered_3_ready =
    xbar_out_3_aw_ready & xbar_awOut_3_io_enq_bits_allowed_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAWOI_filtered_1_3_ready =
    xbar_out_3_aw_ready & xbar_awOut_3_io_enq_bits_allowed_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_3_aw_valid =
    xbar_awOut_3_io_enq_bits_idle
      ? xbar_awOut_3_io_enq_bits_anyValid
      : xbar_awOut_3_io_enq_bits_state_0 & xbar_portsAWOI_filtered_3_valid
        | xbar_awOut_3_io_enq_bits_state_1 & xbar_portsAWOI_filtered_1_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_qos =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_qos : 4'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_3_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_prot =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_prot : 3'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_3_bits_prot
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_cache =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_cache : 4'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_3_bits_cache
         : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_lock =
    xbar_awOut_3_io_enq_bits_muxState_0 & xbar_portsAWOI_filtered_3_bits_lock
    | xbar_awOut_3_io_enq_bits_muxState_1 & xbar_portsAWOI_filtered_1_3_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_burst =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_burst : 2'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_3_bits_burst
         : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_size =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_size : 3'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_3_bits_size
         : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_len =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_len : 8'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_3_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_addr =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_addr : 30'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1
         ? xbar_portsAWOI_filtered_1_3_bits_addr
         : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_aw_bits_id =
    (xbar_awOut_3_io_enq_bits_muxState_0 ? xbar_portsAWOI_filtered_3_bits_id : 3'h0)
    | (xbar_awOut_3_io_enq_bits_muxState_1 ? xbar_portsAWOI_filtered_1_3_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_awOut_3_io_enq_bits =
    {xbar_awOut_3_io_enq_bits_muxState_1, xbar_awOut_3_io_enq_bits_muxState_0};	// src/main/scala/amba/axi4/Xbar.scala:213:81, :292:23
  reg          xbar_idle_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid_3 =
    xbar_portsAROI_filtered_3_valid | xbar_portsAROI_filtered_1_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_valid_3 =
    {xbar_portsAROI_filtered_1_3_valid, xbar_portsAROI_filtered_3_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [1:0]   xbar_readys_mask_3;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [3:0]   xbar_readys_filter_3 =
    {xbar_readys_valid_3 & ~xbar_readys_mask_3, xbar_readys_valid_3};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [3:0]   xbar_readys_unready_3 =
    {xbar_readys_mask_3[1],
     xbar_readys_filter_3[3] | xbar_readys_mask_3[0],
     xbar_readys_filter_3[2:1] | xbar_readys_filter_3[3:2]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:{43,48}
  wire [1:0]   xbar_readys_readys_3 =
    ~(xbar_readys_unready_3[3:2] & xbar_readys_unready_3[1:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_3_0 = xbar_readys_readys_3[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_3_1 = xbar_readys_readys_3[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_3_0 = xbar_readys_3_0 & xbar_portsAROI_filtered_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_3_1 = xbar_readys_3_1 & xbar_portsAROI_filtered_1_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1_3 = xbar_winner_3_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_state_3_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_3_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_3_0 = xbar_idle_3 ? xbar_winner_3_0 : xbar_state_3_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_3_1 = xbar_idle_3 ? xbar_winner_3_1 : xbar_state_3_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_3_0 = xbar_idle_3 ? xbar_readys_3_0 : xbar_state_3_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_3_1 = xbar_idle_3 ? xbar_readys_3_1 : xbar_state_3_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsAROI_filtered_3_ready = xbar_out_3_ar_ready & xbar_allowed_3_0;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_portsAROI_filtered_1_3_ready = xbar_out_3_ar_ready & xbar_allowed_3_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :300:24, :302:31
  assign xbar_out_3_ar_valid =
    xbar_idle_3
      ? xbar_anyValid_3
      : xbar_state_3_0 & xbar_portsAROI_filtered_3_valid | xbar_state_3_1
        & xbar_portsAROI_filtered_1_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_qos =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_qos : 4'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_qos : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_prot =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_prot : 3'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_prot : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_cache =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_cache : 4'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_cache : 4'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_lock =
    xbar_muxState_3_0 & xbar_portsAROI_filtered_3_bits_lock | xbar_muxState_3_1
    & xbar_portsAROI_filtered_1_3_bits_lock;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_burst =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_burst : 2'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_burst : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_size =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_size : 3'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_size : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_len =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_len : 8'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_len : 8'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_addr =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_addr : 30'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_addr : 30'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_ar_bits_id =
    (xbar_muxState_3_0 ? xbar_portsAROI_filtered_3_bits_id : 3'h0)
    | (xbar_muxState_3_1 ? xbar_portsAROI_filtered_1_3_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_out_3_w_valid =
    xbar_awOut_3_io_deq_bits[0] & xbar_portsWOI_filtered_3_valid
    | xbar_awOut_3_io_deq_bits[1] & xbar_portsWOI_filtered_1_3_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_3_w_bits_last =
    xbar_awOut_3_io_deq_bits[0] & xbar_portsWOI_filtered_3_bits_last
    | xbar_awOut_3_io_deq_bits[1] & xbar_portsWOI_filtered_1_3_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_3_w_bits_strb =
    (xbar_awOut_3_io_deq_bits[0] ? xbar_portsWOI_filtered_3_bits_strb : 16'h0)
    | (xbar_awOut_3_io_deq_bits[1] ? xbar_portsWOI_filtered_1_3_bits_strb : 16'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_out_3_w_bits_data =
    (xbar_awOut_3_io_deq_bits[0] ? xbar_portsWOI_filtered_3_bits_data : 128'h0)
    | (xbar_awOut_3_io_deq_bits[1] ? xbar_portsWOI_filtered_1_3_bits_data : 128'h0);	// src/main/scala/amba/axi4/Xbar.scala:178:19, :249:24, src/main/scala/chisel3/util/Mux.scala:30:73, :32:36
  assign xbar_portsWOI_filtered_3_ready =
    xbar_out_3_w_ready & xbar_awOut_3_io_deq_bits[0];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  assign xbar_portsWOI_filtered_1_3_ready =
    xbar_out_3_w_ready & xbar_awOut_3_io_deq_bits[1];	// src/main/scala/amba/axi4/Xbar.scala:178:19, :220:37, :249:24, src/main/scala/chisel3/util/Mux.scala:32:36
  reg          xbar_idle_4;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid_4 =
    xbar_portsRIO_filtered_0_valid | xbar_portsRIO_filtered_1_0_valid
    | xbar_portsRIO_filtered_2_0_valid | xbar_portsRIO_filtered_3_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_lo =
    {xbar_portsRIO_filtered_1_0_valid, xbar_portsRIO_filtered_0_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [1:0]   xbar_readys_hi =
    {xbar_portsRIO_filtered_3_0_valid, xbar_portsRIO_filtered_2_0_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [3:0]   xbar_readys_valid_4 = {xbar_readys_hi, xbar_readys_lo};	// src/main/scala/amba/axi4/Xbar.scala:278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [3:0]   xbar_readys_mask_4;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [7:0]   xbar_readys_filter_4 =
    {xbar_readys_valid_4 & ~xbar_readys_mask_4, xbar_readys_valid_4};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [5:0]   _GEN_6 = xbar_readys_filter_4[6:1] | xbar_readys_filter_4[7:2];	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [4:0]   _GEN_7 = _GEN_6[4:0] | {xbar_readys_filter_4[7], _GEN_6[5:2]};	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [7:0]   xbar_readys_unready_4 =
    {xbar_readys_mask_4[3],
     xbar_readys_filter_4[7] | xbar_readys_mask_4[2],
     _GEN_6[5] | xbar_readys_mask_4[1],
     _GEN_7[4] | xbar_readys_mask_4[0],
     _GEN_7[3:0]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:43
  wire [3:0]   xbar_readys_readys_4 =
    ~(xbar_readys_unready_4[7:4] & xbar_readys_unready_4[3:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_4_0 = xbar_readys_readys_4[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_4_1 = xbar_readys_readys_4[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_4_2 = xbar_readys_readys_4[2];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_4_3 = xbar_readys_readys_4[3];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_4_0 = xbar_readys_4_0 & xbar_portsRIO_filtered_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_4_1 = xbar_readys_4_1 & xbar_portsRIO_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_4_2 = xbar_readys_4_2 & xbar_portsRIO_filtered_2_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_4_3 = xbar_readys_4_3 & xbar_portsRIO_filtered_3_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1_4 = xbar_winner_4_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_2 = xbar_prefixOR_1_4 | xbar_winner_4_1;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_3 = xbar_prefixOR_2 | xbar_winner_4_2;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_state_4_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_4_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_4_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_4_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_4_0 = xbar_idle_4 ? xbar_winner_4_0 : xbar_state_4_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_4_1 = xbar_idle_4 ? xbar_winner_4_1 : xbar_state_4_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_4_2 = xbar_idle_4 ? xbar_winner_4_2 : xbar_state_4_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_4_3 = xbar_idle_4 ? xbar_winner_4_3 : xbar_state_4_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_4_0 = xbar_idle_4 ? xbar_readys_4_0 : xbar_state_4_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_4_1 = xbar_idle_4 ? xbar_readys_4_1 : xbar_state_4_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_4_2 = xbar_idle_4 ? xbar_readys_4_2 : xbar_state_4_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_4_3 = xbar_idle_4 ? xbar_readys_4_3 : xbar_state_4_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsRIO_filtered_0_ready = xbar_in_0_r_ready & xbar_allowed_4_0;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsRIO_filtered_1_0_ready = xbar_in_0_r_ready & xbar_allowed_4_1;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsRIO_filtered_2_0_ready = xbar_in_0_r_ready & xbar_allowed_4_2;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsRIO_filtered_3_0_ready = xbar_in_0_r_ready & xbar_allowed_4_3;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_in_0_r_valid =
    xbar_idle_4
      ? xbar_anyValid_4
      : xbar_state_4_0 & xbar_portsRIO_filtered_0_valid | xbar_state_4_1
        & xbar_portsRIO_filtered_1_0_valid | xbar_state_4_2
        & xbar_portsRIO_filtered_2_0_valid | xbar_state_4_3
        & xbar_portsRIO_filtered_3_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_0_r_bits_last =
    xbar_muxState_4_0 & xbar_portsRIO_filtered_0_bits_last | xbar_muxState_4_1
    & xbar_portsRIO_filtered_1_0_bits_last | xbar_muxState_4_2
    & xbar_portsRIO_filtered_2_0_bits_last | xbar_muxState_4_3
    & xbar_portsRIO_filtered_3_0_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_0_r_bits_resp =
    (xbar_muxState_4_0 ? xbar_portsRIO_filtered_0_bits_resp : 2'h0)
    | (xbar_muxState_4_1 ? xbar_portsRIO_filtered_1_0_bits_resp : 2'h0)
    | (xbar_muxState_4_2 ? xbar_portsRIO_filtered_2_0_bits_resp : 2'h0)
    | (xbar_muxState_4_3 ? xbar_portsRIO_filtered_3_0_bits_resp : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_0_r_bits_data =
    (xbar_muxState_4_0 ? xbar_portsRIO_filtered_0_bits_data : 128'h0)
    | (xbar_muxState_4_1 ? xbar_portsRIO_filtered_1_0_bits_data : 128'h0)
    | (xbar_muxState_4_2 ? xbar_portsRIO_filtered_2_0_bits_data : 128'h0)
    | (xbar_muxState_4_3 ? xbar_portsRIO_filtered_3_0_bits_data : 128'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  wire [2:0]   xbar_in_0_r_bits_id =
    (xbar_muxState_4_0 ? xbar_portsRIO_filtered_0_bits_id : 3'h0)
    | (xbar_muxState_4_1 ? xbar_portsRIO_filtered_1_0_bits_id : 3'h0)
    | (xbar_muxState_4_2 ? xbar_portsRIO_filtered_2_0_bits_id : 3'h0)
    | (xbar_muxState_4_3 ? xbar_portsRIO_filtered_3_0_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  reg          xbar_idle_5;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid_5 =
    xbar_portsBIO_filtered_0_valid | xbar_portsBIO_filtered_1_0_valid
    | xbar_portsBIO_filtered_2_0_valid | xbar_portsBIO_filtered_3_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_lo_1 =
    {xbar_portsBIO_filtered_1_0_valid, xbar_portsBIO_filtered_0_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [1:0]   xbar_readys_hi_1 =
    {xbar_portsBIO_filtered_3_0_valid, xbar_portsBIO_filtered_2_0_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [3:0]   xbar_readys_valid_5 = {xbar_readys_hi_1, xbar_readys_lo_1};	// src/main/scala/amba/axi4/Xbar.scala:278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [3:0]   xbar_readys_mask_5;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [7:0]   xbar_readys_filter_5 =
    {xbar_readys_valid_5 & ~xbar_readys_mask_5, xbar_readys_valid_5};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [5:0]   _GEN_8 = xbar_readys_filter_5[6:1] | xbar_readys_filter_5[7:2];	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [4:0]   _GEN_9 = _GEN_8[4:0] | {xbar_readys_filter_5[7], _GEN_8[5:2]};	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [7:0]   xbar_readys_unready_5 =
    {xbar_readys_mask_5[3],
     xbar_readys_filter_5[7] | xbar_readys_mask_5[2],
     _GEN_8[5] | xbar_readys_mask_5[1],
     _GEN_9[4] | xbar_readys_mask_5[0],
     _GEN_9[3:0]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:43
  wire [3:0]   xbar_readys_readys_5 =
    ~(xbar_readys_unready_5[7:4] & xbar_readys_unready_5[3:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_5_0 = xbar_readys_readys_5[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_5_1 = xbar_readys_readys_5[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_5_2 = xbar_readys_readys_5[2];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_5_3 = xbar_readys_readys_5[3];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_5_0 = xbar_readys_5_0 & xbar_portsBIO_filtered_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_5_1 = xbar_readys_5_1 & xbar_portsBIO_filtered_1_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_5_2 = xbar_readys_5_2 & xbar_portsBIO_filtered_2_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_5_3 = xbar_readys_5_3 & xbar_portsBIO_filtered_3_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1_5 = xbar_winner_5_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_2_1 = xbar_prefixOR_1_5 | xbar_winner_5_1;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_3_1 = xbar_prefixOR_2_1 | xbar_winner_5_2;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_state_5_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_5_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_5_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_5_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_5_0 = xbar_idle_5 ? xbar_winner_5_0 : xbar_state_5_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_5_1 = xbar_idle_5 ? xbar_winner_5_1 : xbar_state_5_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_5_2 = xbar_idle_5 ? xbar_winner_5_2 : xbar_state_5_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_5_3 = xbar_idle_5 ? xbar_winner_5_3 : xbar_state_5_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_5_0 = xbar_idle_5 ? xbar_readys_5_0 : xbar_state_5_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_5_1 = xbar_idle_5 ? xbar_readys_5_1 : xbar_state_5_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_5_2 = xbar_idle_5 ? xbar_readys_5_2 : xbar_state_5_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_5_3 = xbar_idle_5 ? xbar_readys_5_3 : xbar_state_5_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsBIO_filtered_0_ready = xbar_in_0_b_ready & xbar_allowed_5_0;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsBIO_filtered_1_0_ready = xbar_in_0_b_ready & xbar_allowed_5_1;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsBIO_filtered_2_0_ready = xbar_in_0_b_ready & xbar_allowed_5_2;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsBIO_filtered_3_0_ready = xbar_in_0_b_ready & xbar_allowed_5_3;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_in_0_b_valid =
    xbar_idle_5
      ? xbar_anyValid_5
      : xbar_state_5_0 & xbar_portsBIO_filtered_0_valid | xbar_state_5_1
        & xbar_portsBIO_filtered_1_0_valid | xbar_state_5_2
        & xbar_portsBIO_filtered_2_0_valid | xbar_state_5_3
        & xbar_portsBIO_filtered_3_0_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_0_b_bits_resp =
    (xbar_muxState_5_0 ? xbar_portsBIO_filtered_0_bits_resp : 2'h0)
    | (xbar_muxState_5_1 ? xbar_portsBIO_filtered_1_0_bits_resp : 2'h0)
    | (xbar_muxState_5_2 ? xbar_portsBIO_filtered_2_0_bits_resp : 2'h0)
    | (xbar_muxState_5_3 ? xbar_portsBIO_filtered_3_0_bits_resp : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  wire [2:0]   xbar_in_0_b_bits_id =
    (xbar_muxState_5_0 ? xbar_portsBIO_filtered_0_bits_id : 3'h0)
    | (xbar_muxState_5_1 ? xbar_portsBIO_filtered_1_0_bits_id : 3'h0)
    | (xbar_muxState_5_2 ? xbar_portsBIO_filtered_2_0_bits_id : 3'h0)
    | (xbar_muxState_5_3 ? xbar_portsBIO_filtered_3_0_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  reg          xbar_idle_6;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid_6 =
    xbar_portsRIO_filtered_1_valid | xbar_portsRIO_filtered_1_1_valid
    | xbar_portsRIO_filtered_2_1_valid | xbar_portsRIO_filtered_3_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_lo_2 =
    {xbar_portsRIO_filtered_1_1_valid, xbar_portsRIO_filtered_1_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [1:0]   xbar_readys_hi_2 =
    {xbar_portsRIO_filtered_3_1_valid, xbar_portsRIO_filtered_2_1_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [3:0]   xbar_readys_valid_6 = {xbar_readys_hi_2, xbar_readys_lo_2};	// src/main/scala/amba/axi4/Xbar.scala:278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [3:0]   xbar_readys_mask_6;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [7:0]   xbar_readys_filter_6 =
    {xbar_readys_valid_6 & ~xbar_readys_mask_6, xbar_readys_valid_6};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [5:0]   _GEN_10 = xbar_readys_filter_6[6:1] | xbar_readys_filter_6[7:2];	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [4:0]   _GEN_11 = _GEN_10[4:0] | {xbar_readys_filter_6[7], _GEN_10[5:2]};	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [7:0]   xbar_readys_unready_6 =
    {xbar_readys_mask_6[3],
     xbar_readys_filter_6[7] | xbar_readys_mask_6[2],
     _GEN_10[5] | xbar_readys_mask_6[1],
     _GEN_11[4] | xbar_readys_mask_6[0],
     _GEN_11[3:0]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:43
  wire [3:0]   xbar_readys_readys_6 =
    ~(xbar_readys_unready_6[7:4] & xbar_readys_unready_6[3:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_6_0 = xbar_readys_readys_6[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_6_1 = xbar_readys_readys_6[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_6_2 = xbar_readys_readys_6[2];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_6_3 = xbar_readys_readys_6[3];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_6_0 = xbar_readys_6_0 & xbar_portsRIO_filtered_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_6_1 = xbar_readys_6_1 & xbar_portsRIO_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_6_2 = xbar_readys_6_2 & xbar_portsRIO_filtered_2_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_6_3 = xbar_readys_6_3 & xbar_portsRIO_filtered_3_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1_6 = xbar_winner_6_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_2_2 = xbar_prefixOR_1_6 | xbar_winner_6_1;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_3_2 = xbar_prefixOR_2_2 | xbar_winner_6_2;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  reg          xbar_state_6_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_6_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_6_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_6_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_6_0 = xbar_idle_6 ? xbar_winner_6_0 : xbar_state_6_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_6_1 = xbar_idle_6 ? xbar_winner_6_1 : xbar_state_6_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_6_2 = xbar_idle_6 ? xbar_winner_6_2 : xbar_state_6_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_6_3 = xbar_idle_6 ? xbar_winner_6_3 : xbar_state_6_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_6_0 = xbar_idle_6 ? xbar_readys_6_0 : xbar_state_6_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_6_1 = xbar_idle_6 ? xbar_readys_6_1 : xbar_state_6_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_6_2 = xbar_idle_6 ? xbar_readys_6_2 : xbar_state_6_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_6_3 = xbar_idle_6 ? xbar_readys_6_3 : xbar_state_6_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsRIO_filtered_1_ready = xbar_in_1_r_ready & xbar_allowed_6_0;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsRIO_filtered_1_1_ready = xbar_in_1_r_ready & xbar_allowed_6_1;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsRIO_filtered_2_1_ready = xbar_in_1_r_ready & xbar_allowed_6_2;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsRIO_filtered_3_1_ready = xbar_in_1_r_ready & xbar_allowed_6_3;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_in_1_r_valid =
    xbar_idle_6
      ? xbar_anyValid_6
      : xbar_state_6_0 & xbar_portsRIO_filtered_1_valid | xbar_state_6_1
        & xbar_portsRIO_filtered_1_1_valid | xbar_state_6_2
        & xbar_portsRIO_filtered_2_1_valid | xbar_state_6_3
        & xbar_portsRIO_filtered_3_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_1_r_bits_last =
    xbar_muxState_6_0 & xbar_portsRIO_filtered_1_bits_last | xbar_muxState_6_1
    & xbar_portsRIO_filtered_1_1_bits_last | xbar_muxState_6_2
    & xbar_portsRIO_filtered_2_1_bits_last | xbar_muxState_6_3
    & xbar_portsRIO_filtered_3_1_bits_last;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_1_r_bits_resp =
    (xbar_muxState_6_0 ? xbar_portsRIO_filtered_1_bits_resp : 2'h0)
    | (xbar_muxState_6_1 ? xbar_portsRIO_filtered_1_1_bits_resp : 2'h0)
    | (xbar_muxState_6_2 ? xbar_portsRIO_filtered_2_1_bits_resp : 2'h0)
    | (xbar_muxState_6_3 ? xbar_portsRIO_filtered_3_1_bits_resp : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_1_r_bits_data =
    (xbar_muxState_6_0 ? xbar_portsRIO_filtered_1_bits_data : 128'h0)
    | (xbar_muxState_6_1 ? xbar_portsRIO_filtered_1_1_bits_data : 128'h0)
    | (xbar_muxState_6_2 ? xbar_portsRIO_filtered_2_1_bits_data : 128'h0)
    | (xbar_muxState_6_3 ? xbar_portsRIO_filtered_3_1_bits_data : 128'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_1_r_bits_id =
    (xbar_muxState_6_0 ? xbar_portsRIO_filtered_1_bits_id : 3'h0)
    | (xbar_muxState_6_1 ? xbar_portsRIO_filtered_1_1_bits_id : 3'h0)
    | (xbar_muxState_6_2 ? xbar_portsRIO_filtered_2_1_bits_id : 3'h0)
    | (xbar_muxState_6_3 ? xbar_portsRIO_filtered_3_1_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  reg          xbar_idle_7;	// src/main/scala/amba/axi4/Xbar.scala:272:23
  wire         xbar_anyValid_7 =
    xbar_portsBIO_filtered_1_valid | xbar_portsBIO_filtered_1_1_valid
    | xbar_portsBIO_filtered_2_1_valid | xbar_portsBIO_filtered_3_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :276:36
  wire [1:0]   xbar_readys_lo_3 =
    {xbar_portsBIO_filtered_1_1_valid, xbar_portsBIO_filtered_1_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [1:0]   xbar_readys_hi_3 =
    {xbar_portsBIO_filtered_3_1_valid, xbar_portsBIO_filtered_2_1_valid};	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:49
  wire [3:0]   xbar_readys_valid_7 = {xbar_readys_hi_3, xbar_readys_lo_3};	// src/main/scala/amba/axi4/Xbar.scala:278:49, src/main/scala/tilelink/Arbiter.scala:21:23
  reg  [3:0]   xbar_readys_mask_7;	// src/main/scala/tilelink/Arbiter.scala:23:23
  wire [7:0]   xbar_readys_filter_7 =
    {xbar_readys_valid_7 & ~xbar_readys_mask_7, xbar_readys_valid_7};	// src/main/scala/tilelink/Arbiter.scala:21:23, :23:23, :24:{21,28,30}
  wire [5:0]   _GEN_12 = xbar_readys_filter_7[6:1] | xbar_readys_filter_7[7:2];	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [4:0]   _GEN_13 = _GEN_12[4:0] | {xbar_readys_filter_7[7], _GEN_12[5:2]};	// src/main/scala/tilelink/Arbiter.scala:24:21, src/main/scala/util/package.scala:262:{43,48}
  wire [7:0]   xbar_readys_unready_7 =
    {xbar_readys_mask_7[3],
     xbar_readys_filter_7[7] | xbar_readys_mask_7[2],
     _GEN_12[5] | xbar_readys_mask_7[1],
     _GEN_13[4] | xbar_readys_mask_7[0],
     _GEN_13[3:0]};	// src/main/scala/tilelink/Arbiter.scala:23:23, :24:21, :25:58, src/main/scala/util/package.scala:262:43
  wire [3:0]   xbar_readys_readys_7 =
    ~(xbar_readys_unready_7[7:4] & xbar_readys_unready_7[3:0]);	// src/main/scala/tilelink/Arbiter.scala:25:58, :26:{18,29,39,48}
  wire         xbar_readys_7_0 = xbar_readys_readys_7[0];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_7_1 = xbar_readys_readys_7[1];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_7_2 = xbar_readys_readys_7[2];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_readys_7_3 = xbar_readys_readys_7[3];	// src/main/scala/amba/axi4/Xbar.scala:278:{25,73}, src/main/scala/tilelink/Arbiter.scala:26:18
  wire         xbar_winner_7_0 = xbar_readys_7_0 & xbar_portsBIO_filtered_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_7_1 = xbar_readys_7_1 & xbar_portsBIO_filtered_1_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_7_2 = xbar_readys_7_2 & xbar_portsBIO_filtered_2_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_winner_7_3 = xbar_readys_7_3 & xbar_portsBIO_filtered_3_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:249:24, :278:25, :280:{25,67}
  wire         xbar_prefixOR_1_7 = xbar_winner_7_0;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_2_3 = xbar_prefixOR_1_7 | xbar_winner_7_1;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  wire         xbar_prefixOR_3_3 = xbar_prefixOR_2_3 | xbar_winner_7_2;	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46
  `ifndef SYNTHESIS	// src/main/scala/amba/axi4/Xbar.scala:131:22
    always @(posedge clock) begin	// src/main/scala/amba/axi4/Xbar.scala:131:22
      if (~reset & ~(~xbar__arFIFOMap_0_T_4 | (|xbar_arFIFOMap_0_count))) begin	// src/main/scala/amba/axi4/Xbar.scala:128:34, :131:{22,23,34,43}, :144:43, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $error("Assertion failed\n    at Xbar.scala:131 assert (!resp_fire || count =/= 0.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:131:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:131:22
      end
      if (~reset & ~(~xbar__arFIFOMap_0_T | xbar__arFIFOMap_0_T_12)) begin	// src/main/scala/amba/axi4/Xbar.scala:132:{22,23,34,43}, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $error("Assertion failed\n    at Xbar.scala:132 assert (!req_fire  || count =/= flight.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:132:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:132:22
      end
      if (~reset & ~(~xbar__awFIFOMap_0_T_2 | (|xbar_awFIFOMap_0_count))) begin	// src/main/scala/amba/axi4/Xbar.scala:128:34, :131:{22,23,34,43}, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $error("Assertion failed\n    at Xbar.scala:131 assert (!resp_fire || count =/= 0.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:131:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:131:22
      end
      if (~reset & ~(~xbar__awFIFOMap_0_T | xbar__awFIFOMap_0_T_11)) begin	// src/main/scala/amba/axi4/Xbar.scala:132:{22,23,34,43}, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $error("Assertion failed\n    at Xbar.scala:132 assert (!req_fire  || count =/= flight.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:132:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:132:22
      end
      if (~reset & ~(~xbar__arFIFOMap_2_T_6 | (|xbar_arFIFOMap_2_count))) begin	// src/main/scala/amba/axi4/Xbar.scala:128:34, :131:{22,23,34,43}, :144:{24,43}, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $error("Assertion failed\n    at Xbar.scala:131 assert (!resp_fire || count =/= 0.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:131:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:131:22
      end
      if (~reset & ~(~xbar__arFIFOMap_2_T_2 | xbar__arFIFOMap_2_T_14)) begin	// src/main/scala/amba/axi4/Xbar.scala:132:{22,23,34,43}, :143:25, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $error("Assertion failed\n    at Xbar.scala:132 assert (!req_fire  || count =/= flight.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:132:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:132:22
      end
      if (~reset & ~(~xbar__awFIFOMap_2_T_5 | (|xbar_awFIFOMap_2_count))) begin	// src/main/scala/amba/axi4/Xbar.scala:128:34, :131:{22,23,34,43}, :148:24, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $error("Assertion failed\n    at Xbar.scala:131 assert (!resp_fire || count =/= 0.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:131:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:131:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:131:22
      end
      if (~reset & ~(~xbar__awFIFOMap_2_T_2 | xbar__awFIFOMap_2_T_13)) begin	// src/main/scala/amba/axi4/Xbar.scala:132:{22,23,34,43}, :147:25, src/main/scala/chisel3/util/Decoupled.scala:52:35
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $error("Assertion failed\n    at Xbar.scala:132 assert (!req_fire  || count =/= flight.U)\n");	// src/main/scala/amba/axi4/Xbar.scala:132:22
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:132:22
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:132:22
      end
      if (~reset
          & xbar_awOut_0_io_enq_bits_readys_valid != xbar_awOut_0_io_enq_bits_readys_valid) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~(~xbar_awOut_0_io_enq_bits_prefixOR_1
              | ~xbar_awOut_0_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_awOut_0_io_enq_bits_anyValid | xbar_awOut_0_io_enq_bits_winner_0
              | xbar_awOut_0_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid != xbar_readys_valid) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset & ~(~xbar_prefixOR_1 | ~xbar_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset & ~(~xbar_anyValid | xbar_winner_0 | xbar_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset
          & xbar_awOut_1_io_enq_bits_readys_valid != xbar_awOut_1_io_enq_bits_readys_valid) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~(~xbar_awOut_1_io_enq_bits_prefixOR_1
              | ~xbar_awOut_1_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_awOut_1_io_enq_bits_anyValid | xbar_awOut_1_io_enq_bits_winner_0
              | xbar_awOut_1_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid_1 != xbar_readys_valid_1) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset & ~(~xbar_prefixOR_1_1 | ~xbar_winner_1_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset & ~(~xbar_anyValid_1 | xbar_winner_1_0 | xbar_winner_1_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset
          & xbar_awOut_2_io_enq_bits_readys_valid != xbar_awOut_2_io_enq_bits_readys_valid) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~(~xbar_awOut_2_io_enq_bits_prefixOR_1
              | ~xbar_awOut_2_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_awOut_2_io_enq_bits_anyValid | xbar_awOut_2_io_enq_bits_winner_0
              | xbar_awOut_2_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid_2 != xbar_readys_valid_2) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset & ~(~xbar_prefixOR_1_2 | ~xbar_winner_2_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset & ~(~xbar_anyValid_2 | xbar_winner_2_0 | xbar_winner_2_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset
          & xbar_awOut_3_io_enq_bits_readys_valid != xbar_awOut_3_io_enq_bits_readys_valid) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~(~xbar_awOut_3_io_enq_bits_prefixOR_1
              | ~xbar_awOut_3_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_awOut_3_io_enq_bits_anyValid | xbar_awOut_3_io_enq_bits_winner_0
              | xbar_awOut_3_io_enq_bits_winner_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid_3 != xbar_readys_valid_3) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset & ~(~xbar_prefixOR_1_3 | ~xbar_winner_3_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset & ~(~xbar_anyValid_3 | xbar_winner_3_0 | xbar_winner_3_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid_4 != xbar_readys_valid_4) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~((~xbar_prefixOR_1_4 | ~xbar_winner_4_1)
              & (~xbar_prefixOR_2 | ~xbar_winner_4_2)
              & (~xbar_prefixOR_3 | ~xbar_winner_4_3))) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60,75}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_anyValid_4 | xbar_winner_4_0 | xbar_winner_4_1 | xbar_winner_4_2
              | xbar_winner_4_3)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid_5 != xbar_readys_valid_5) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~((~xbar_prefixOR_1_5 | ~xbar_winner_5_1)
              & (~xbar_prefixOR_2_1 | ~xbar_winner_5_2)
              & (~xbar_prefixOR_3_1 | ~xbar_winner_5_3))) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60,75}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_anyValid_5 | xbar_winner_5_0 | xbar_winner_5_1 | xbar_winner_5_2
              | xbar_winner_5_3)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid_6 != xbar_readys_valid_6) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~((~xbar_prefixOR_1_6 | ~xbar_winner_6_1)
              & (~xbar_prefixOR_2_2 | ~xbar_winner_6_2)
              & (~xbar_prefixOR_3_2 | ~xbar_winner_6_3))) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60,75}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_anyValid_6 | xbar_winner_6_0 | xbar_winner_6_1 | xbar_winner_6_2
              | xbar_winner_6_3)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
      if (~reset & xbar_readys_valid_7 != xbar_readys_valid_7) begin	// src/main/scala/tilelink/Arbiter.scala:21:23, :22:{12,19}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");	// src/main/scala/tilelink/Arbiter.scala:22:12
        if (`STOP_COND_)	// src/main/scala/tilelink/Arbiter.scala:22:12
          $fatal;	// src/main/scala/tilelink/Arbiter.scala:22:12
      end
      if (~reset
          & ~((~xbar_prefixOR_1_7 | ~xbar_winner_7_1)
              & (~xbar_prefixOR_2_3 | ~xbar_winner_7_2)
              & (~xbar_prefixOR_3_3 | ~xbar_winner_7_3))) begin	// src/main/scala/amba/axi4/Xbar.scala:280:25, :285:46, :286:{11,54,57,60,75}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $error("Assertion failed\n    at Xbar.scala:286 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");	// src/main/scala/amba/axi4/Xbar.scala:286:11
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:286:11
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:286:11
      end
      if (~reset
          & ~(~xbar_anyValid_7 | xbar_winner_7_0 | xbar_winner_7_1 | xbar_winner_7_2
              | xbar_winner_7_3)) begin	// src/main/scala/amba/axi4/Xbar.scala:276:36, :280:25, :286:11, :288:{12,13,23,41}
        if (`ASSERT_VERBOSE_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $error("Assertion failed\n    at Xbar.scala:288 assert (!anyValid || winner.reduce(_||_))\n");	// src/main/scala/amba/axi4/Xbar.scala:288:12
        if (`STOP_COND_)	// src/main/scala/amba/axi4/Xbar.scala:288:12
          $fatal;	// src/main/scala/amba/axi4/Xbar.scala:288:12
      end
    end // always @(posedge)
  `endif // not def SYNTHESIS
  reg          xbar_state_7_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_7_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_7_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  reg          xbar_state_7_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24
  wire         xbar_muxState_7_0 = xbar_idle_7 ? xbar_winner_7_0 : xbar_state_7_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_7_1 = xbar_idle_7 ? xbar_winner_7_1 : xbar_state_7_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_7_2 = xbar_idle_7 ? xbar_winner_7_2 : xbar_state_7_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_muxState_7_3 = xbar_idle_7 ? xbar_winner_7_3 : xbar_state_7_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :280:25, :291:24, :292:23
  wire         xbar_allowed_7_0 = xbar_idle_7 ? xbar_readys_7_0 : xbar_state_7_0;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_7_1 = xbar_idle_7 ? xbar_readys_7_1 : xbar_state_7_1;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_7_2 = xbar_idle_7 ? xbar_readys_7_2 : xbar_state_7_2;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  wire         xbar_allowed_7_3 = xbar_idle_7 ? xbar_readys_7_3 : xbar_state_7_3;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :278:25, :291:24, :300:24
  assign xbar_portsBIO_filtered_1_ready = xbar_in_1_b_ready & xbar_allowed_7_0;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsBIO_filtered_1_1_ready = xbar_in_1_b_ready & xbar_allowed_7_1;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsBIO_filtered_2_1_ready = xbar_in_1_b_ready & xbar_allowed_7_2;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_portsBIO_filtered_3_1_ready = xbar_in_1_b_ready & xbar_allowed_7_3;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :300:24, :302:31
  assign xbar_in_1_b_valid =
    xbar_idle_7
      ? xbar_anyValid_7
      : xbar_state_7_0 & xbar_portsBIO_filtered_1_valid | xbar_state_7_1
        & xbar_portsBIO_filtered_1_1_valid | xbar_state_7_2
        & xbar_portsBIO_filtered_2_1_valid | xbar_state_7_3
        & xbar_portsBIO_filtered_3_1_valid;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :272:23, :276:36, :291:24, :308:22, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_1_b_bits_resp =
    (xbar_muxState_7_0 ? xbar_portsBIO_filtered_1_bits_resp : 2'h0)
    | (xbar_muxState_7_1 ? xbar_portsBIO_filtered_1_1_bits_resp : 2'h0)
    | (xbar_muxState_7_2 ? xbar_portsBIO_filtered_2_1_bits_resp : 2'h0)
    | (xbar_muxState_7_3 ? xbar_portsBIO_filtered_3_1_bits_resp : 2'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  assign xbar_in_1_b_bits_id =
    (xbar_muxState_7_0 ? xbar_portsBIO_filtered_1_bits_id : 3'h0)
    | (xbar_muxState_7_1 ? xbar_portsBIO_filtered_1_1_bits_id : 3'h0)
    | (xbar_muxState_7_2 ? xbar_portsBIO_filtered_2_1_bits_id : 3'h0)
    | (xbar_muxState_7_3 ? xbar_portsBIO_filtered_3_1_bits_id : 3'h0);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :249:24, :292:23, src/main/scala/chisel3/util/Mux.scala:30:73
  wire         master1_aw_ready_0 = mapMasterOut_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_valid = mapMasterOut_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_id = mapMasterOut_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_addr = mapMasterOut_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_len = mapMasterOut_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_size = mapMasterOut_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_burst = mapMasterOut_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_lock = mapMasterOut_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_cache = mapMasterOut_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_prot = mapMasterOut_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_aw_bits_qos = mapMasterOut_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master1_w_ready_0 = mapMasterOut_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_w_valid = mapMasterOut_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_w_bits_data = mapMasterOut_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_w_bits_strb = mapMasterOut_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_w_bits_last = mapMasterOut_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_b_ready = mapMasterOut_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master1_b_valid_0 = mapMasterOut_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   master1_b_bits_resp_0 = mapMasterOut_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master1_ar_ready_0 = mapMasterOut_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_valid = mapMasterOut_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_id = mapMasterOut_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_addr = mapMasterOut_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_len = mapMasterOut_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_size = mapMasterOut_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_burst = mapMasterOut_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_lock = mapMasterOut_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_cache = mapMasterOut_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_prot = mapMasterOut_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_ar_bits_qos = mapMasterOut_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_0_r_ready = mapMasterOut_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master1_r_valid_0 = mapMasterOut_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] master1_r_bits_data_0 = mapMasterOut_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   master1_r_bits_resp_0 = mapMasterOut_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master1_r_bits_last_0 = mapMasterOut_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master2_aw_ready_0 = mapMasterOut_1_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_valid = mapMasterOut_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_id = mapMasterOut_1_aw_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_addr = mapMasterOut_1_aw_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_len = mapMasterOut_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_size = mapMasterOut_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_burst = mapMasterOut_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_lock = mapMasterOut_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_cache = mapMasterOut_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_prot = mapMasterOut_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_aw_bits_qos = mapMasterOut_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master2_w_ready_0 = mapMasterOut_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_w_valid = mapMasterOut_1_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_w_bits_data = mapMasterOut_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_w_bits_strb = mapMasterOut_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_w_bits_last = mapMasterOut_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_b_ready = mapMasterOut_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master2_b_valid_0 = mapMasterOut_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   master2_b_bits_resp_0 = mapMasterOut_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master2_ar_ready_0 = mapMasterOut_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_valid = mapMasterOut_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_id = mapMasterOut_1_ar_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_addr = mapMasterOut_1_ar_bits_addr;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_len = mapMasterOut_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_size = mapMasterOut_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_burst = mapMasterOut_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_lock = mapMasterOut_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_cache = mapMasterOut_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_prot = mapMasterOut_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_ar_bits_qos = mapMasterOut_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_in_1_r_ready = mapMasterOut_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master2_r_valid_0 = mapMasterOut_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [127:0] master2_r_bits_data_0 = mapMasterOut_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire [1:0]   master2_r_bits_resp_0 = mapMasterOut_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  wire         master2_r_bits_last_0 = mapMasterOut_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17
  assign xbar_auto_anon_out_0_aw_ready = mapSlaveIn_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_aw_valid_0 = mapSlaveIn_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave1_aw_bits_len_0 = mapSlaveIn_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave1_aw_bits_size_0 = mapSlaveIn_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave1_aw_bits_burst_0 = mapSlaveIn_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_aw_bits_lock_0 = mapSlaveIn_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave1_aw_bits_cache_0 = mapSlaveIn_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave1_aw_bits_prot_0 = mapSlaveIn_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave1_aw_bits_qos_0 = mapSlaveIn_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_w_ready = mapSlaveIn_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_w_valid_0 = mapSlaveIn_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] slave1_w_bits_data_0 = mapSlaveIn_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  slave1_w_bits_strb_0 = mapSlaveIn_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_w_bits_last_0 = mapSlaveIn_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_b_ready_0 = mapSlaveIn_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_b_valid = mapSlaveIn_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_b_bits_id = mapSlaveIn_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_b_bits_resp = mapSlaveIn_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_ar_ready = mapSlaveIn_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_ar_valid_0 = mapSlaveIn_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave1_ar_bits_len_0 = mapSlaveIn_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave1_ar_bits_size_0 = mapSlaveIn_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave1_ar_bits_burst_0 = mapSlaveIn_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_ar_bits_lock_0 = mapSlaveIn_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave1_ar_bits_cache_0 = mapSlaveIn_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave1_ar_bits_prot_0 = mapSlaveIn_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave1_ar_bits_qos_0 = mapSlaveIn_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave1_r_ready_0 = mapSlaveIn_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_r_valid = mapSlaveIn_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_r_bits_id = mapSlaveIn_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_r_bits_data = mapSlaveIn_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_r_bits_resp = mapSlaveIn_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_0_r_bits_last = mapSlaveIn_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_aw_ready = mapSlaveIn_1_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_aw_valid_0 = mapSlaveIn_1_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave2_aw_bits_len_0 = mapSlaveIn_1_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave2_aw_bits_size_0 = mapSlaveIn_1_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave2_aw_bits_burst_0 = mapSlaveIn_1_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_aw_bits_lock_0 = mapSlaveIn_1_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave2_aw_bits_cache_0 = mapSlaveIn_1_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave2_aw_bits_prot_0 = mapSlaveIn_1_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave2_aw_bits_qos_0 = mapSlaveIn_1_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_w_ready = mapSlaveIn_1_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_w_valid_0 = mapSlaveIn_1_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] slave2_w_bits_data_0 = mapSlaveIn_1_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  slave2_w_bits_strb_0 = mapSlaveIn_1_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_w_bits_last_0 = mapSlaveIn_1_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_b_ready_0 = mapSlaveIn_1_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_b_valid = mapSlaveIn_1_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_b_bits_id = mapSlaveIn_1_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_b_bits_resp = mapSlaveIn_1_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_ar_ready = mapSlaveIn_1_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_ar_valid_0 = mapSlaveIn_1_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave2_ar_bits_len_0 = mapSlaveIn_1_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave2_ar_bits_size_0 = mapSlaveIn_1_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave2_ar_bits_burst_0 = mapSlaveIn_1_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_ar_bits_lock_0 = mapSlaveIn_1_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave2_ar_bits_cache_0 = mapSlaveIn_1_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave2_ar_bits_prot_0 = mapSlaveIn_1_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave2_ar_bits_qos_0 = mapSlaveIn_1_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave2_r_ready_0 = mapSlaveIn_1_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_r_valid = mapSlaveIn_1_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_r_bits_id = mapSlaveIn_1_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_r_bits_data = mapSlaveIn_1_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_r_bits_resp = mapSlaveIn_1_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_1_r_bits_last = mapSlaveIn_1_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_aw_ready = mapSlaveIn_2_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_aw_valid_0 = mapSlaveIn_2_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave3_aw_bits_len_0 = mapSlaveIn_2_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave3_aw_bits_size_0 = mapSlaveIn_2_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave3_aw_bits_burst_0 = mapSlaveIn_2_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_aw_bits_lock_0 = mapSlaveIn_2_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave3_aw_bits_cache_0 = mapSlaveIn_2_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave3_aw_bits_prot_0 = mapSlaveIn_2_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave3_aw_bits_qos_0 = mapSlaveIn_2_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_w_ready = mapSlaveIn_2_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_w_valid_0 = mapSlaveIn_2_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] slave3_w_bits_data_0 = mapSlaveIn_2_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  slave3_w_bits_strb_0 = mapSlaveIn_2_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_w_bits_last_0 = mapSlaveIn_2_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_b_ready_0 = mapSlaveIn_2_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_b_valid = mapSlaveIn_2_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_b_bits_id = mapSlaveIn_2_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_b_bits_resp = mapSlaveIn_2_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_ar_ready = mapSlaveIn_2_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_ar_valid_0 = mapSlaveIn_2_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave3_ar_bits_len_0 = mapSlaveIn_2_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave3_ar_bits_size_0 = mapSlaveIn_2_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave3_ar_bits_burst_0 = mapSlaveIn_2_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_ar_bits_lock_0 = mapSlaveIn_2_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave3_ar_bits_cache_0 = mapSlaveIn_2_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave3_ar_bits_prot_0 = mapSlaveIn_2_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave3_ar_bits_qos_0 = mapSlaveIn_2_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave3_r_ready_0 = mapSlaveIn_2_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_r_valid = mapSlaveIn_2_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_r_bits_id = mapSlaveIn_2_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_r_bits_data = mapSlaveIn_2_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_r_bits_resp = mapSlaveIn_2_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_2_r_bits_last = mapSlaveIn_2_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_aw_ready = mapSlaveIn_3_aw_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_aw_valid_0 = mapSlaveIn_3_aw_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave4_aw_bits_len_0 = mapSlaveIn_3_aw_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave4_aw_bits_size_0 = mapSlaveIn_3_aw_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave4_aw_bits_burst_0 = mapSlaveIn_3_aw_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_aw_bits_lock_0 = mapSlaveIn_3_aw_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave4_aw_bits_cache_0 = mapSlaveIn_3_aw_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave4_aw_bits_prot_0 = mapSlaveIn_3_aw_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave4_aw_bits_qos_0 = mapSlaveIn_3_aw_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_w_ready = mapSlaveIn_3_w_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_w_valid_0 = mapSlaveIn_3_w_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [127:0] slave4_w_bits_data_0 = mapSlaveIn_3_w_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [15:0]  slave4_w_bits_strb_0 = mapSlaveIn_3_w_bits_strb;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_w_bits_last_0 = mapSlaveIn_3_w_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_b_ready_0 = mapSlaveIn_3_b_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_b_valid = mapSlaveIn_3_b_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_b_bits_id = mapSlaveIn_3_b_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_b_bits_resp = mapSlaveIn_3_b_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_ar_ready = mapSlaveIn_3_ar_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_ar_valid_0 = mapSlaveIn_3_ar_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [7:0]   slave4_ar_bits_len_0 = mapSlaveIn_3_ar_bits_len;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave4_ar_bits_size_0 = mapSlaveIn_3_ar_bits_size;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [1:0]   slave4_ar_bits_burst_0 = mapSlaveIn_3_ar_bits_burst;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_ar_bits_lock_0 = mapSlaveIn_3_ar_bits_lock;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave4_ar_bits_cache_0 = mapSlaveIn_3_ar_bits_cache;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [2:0]   slave4_ar_bits_prot_0 = mapSlaveIn_3_ar_bits_prot;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire [3:0]   slave4_ar_bits_qos_0 = mapSlaveIn_3_ar_bits_qos;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  wire         slave4_r_ready_0 = mapSlaveIn_3_r_ready;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_r_valid = mapSlaveIn_3_r_valid;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_r_bits_id = mapSlaveIn_3_r_bits_id;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_r_bits_data = mapSlaveIn_3_r_bits_data;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_r_bits_resp = mapSlaveIn_3_r_bits_resp;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign xbar_auto_anon_out_3_r_bits_last = mapSlaveIn_3_r_bits_last;	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17
  assign mapMasterOut_aw_bits_id = master1_aw_bits_id_0[0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  assign mapMasterOut_aw_bits_addr = master1_aw_bits_addr_0[29:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  assign mapMasterOut_ar_bits_id = master1_ar_bits_id_0[0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  assign mapMasterOut_ar_bits_addr = master1_ar_bits_addr_0[29:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  assign mapMasterOut_1_aw_bits_id = master2_aw_bits_id_0[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  assign mapMasterOut_1_aw_bits_addr = master2_aw_bits_addr_0[29:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  wire [7:0]   master2_b_bits_id_0 = {6'h0, mapMasterOut_1_b_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  assign mapMasterOut_1_ar_bits_id = master2_ar_bits_id_0[1:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  assign mapMasterOut_1_ar_bits_addr = master2_ar_bits_addr_0[29:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  wire [7:0]   master2_r_bits_id_0 = {6'h0, mapMasterOut_1_r_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:542:17, src/main/scala/componentgen/componentgenModule.scala:72:33
  wire [7:0]   slave1_aw_bits_id_0 = {5'h0, mapSlaveIn_aw_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave1_aw_bits_addr_0 = {20'h0, mapSlaveIn_aw_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_b_bits_id = slave1_b_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [7:0]   slave1_ar_bits_id_0 = {5'h0, mapSlaveIn_ar_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave1_ar_bits_addr_0 = {20'h0, mapSlaveIn_ar_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_r_bits_id = slave1_r_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [7:0]   slave2_aw_bits_id_0 = {5'h0, mapSlaveIn_1_aw_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave2_aw_bits_addr_0 = {19'h0, mapSlaveIn_1_aw_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_1_b_bits_id = slave2_b_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [7:0]   slave2_ar_bits_id_0 = {5'h0, mapSlaveIn_1_ar_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave2_ar_bits_addr_0 = {19'h0, mapSlaveIn_1_ar_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_1_r_bits_id = slave2_r_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [7:0]   slave3_aw_bits_id_0 = {5'h0, mapSlaveIn_2_aw_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave3_aw_bits_addr_0 = {18'h0, mapSlaveIn_2_aw_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_2_b_bits_id = slave3_b_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [7:0]   slave3_ar_bits_id_0 = {5'h0, mapSlaveIn_2_ar_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave3_ar_bits_addr_0 = {18'h0, mapSlaveIn_2_ar_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_2_r_bits_id = slave3_r_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [7:0]   slave4_aw_bits_id_0 = {5'h0, mapSlaveIn_3_aw_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave4_aw_bits_addr_0 = {18'h0, mapSlaveIn_3_aw_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_3_b_bits_id = slave4_b_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [7:0]   slave4_ar_bits_id_0 = {5'h0, mapSlaveIn_3_ar_bits_id};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  wire [47:0]  slave4_ar_bits_addr_0 = {18'h0, mapSlaveIn_3_ar_bits_addr};	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  assign mapSlaveIn_3_r_bits_id = slave4_r_bits_id_0[2:0];	// dependencies/diplomacy/diplomacy/src/diplomacy/nodes/MixedNode.scala:551:17, src/main/scala/componentgen/componentgenModule.scala:77:31
  always @(posedge clock) begin
    if (reset) begin
      xbar_awIn_0_enq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awIn_0_deq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awIn_0_maybe_full <= 1'h0;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
      xbar_awIn_1_enq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awIn_1_deq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awIn_1_maybe_full <= 1'h0;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
      xbar_awOut_0_enq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_0_deq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_0_maybe_full <= 1'h0;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
      xbar_awOut_1_enq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_1_deq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_1_maybe_full <= 1'h0;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
      xbar_awOut_2_enq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_2_deq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_2_maybe_full <= 1'h0;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
      xbar_awOut_3_enq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_3_deq_ptr_value <= 1'h0;	// src/main/scala/chisel3/util/Counter.scala:61:40
      xbar_awOut_3_maybe_full <= 1'h0;	// src/main/scala/chisel3/util/Decoupled.scala:260:27
      xbar_arFIFOMap_0_count <= 3'h0;	// src/main/scala/amba/axi4/Xbar.scala:128:34
      xbar_awFIFOMap_0_count <= 3'h0;	// src/main/scala/amba/axi4/Xbar.scala:128:34
      xbar_latched <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:161:30
      xbar_arFIFOMap_2_count <= 3'h0;	// src/main/scala/amba/axi4/Xbar.scala:128:34
      xbar_awFIFOMap_2_count <= 3'h0;	// src/main/scala/amba/axi4/Xbar.scala:128:34
      xbar_latched_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:161:30
      xbar_latched_2 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:186:30
      xbar_latched_3 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:186:30
      xbar_latched_4 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:186:30
      xbar_latched_5 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:186:30
      xbar_awOut_0_io_enq_bits_idle <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_awOut_0_io_enq_bits_readys_mask <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_awOut_0_io_enq_bits_state_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_awOut_0_io_enq_bits_state_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_awOut_1_io_enq_bits_idle <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_awOut_1_io_enq_bits_readys_mask <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_awOut_1_io_enq_bits_state_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_awOut_1_io_enq_bits_state_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle_1 <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask_1 <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_1_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_1_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_awOut_2_io_enq_bits_idle <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_awOut_2_io_enq_bits_readys_mask <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_awOut_2_io_enq_bits_state_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_awOut_2_io_enq_bits_state_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle_2 <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask_2 <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_2_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_2_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_awOut_3_io_enq_bits_idle <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_awOut_3_io_enq_bits_readys_mask <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_awOut_3_io_enq_bits_state_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_awOut_3_io_enq_bits_state_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle_3 <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask_3 <= 2'h3;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_3_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_3_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle_4 <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask_4 <= 4'hF;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_4_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_4_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_4_2 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_4_3 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle_5 <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask_5 <= 4'hF;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_5_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_5_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_5_2 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_5_3 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle_6 <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask_6 <= 4'hF;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_6_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_6_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_6_2 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_6_3 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_idle_7 <= 1'h1;	// src/main/scala/amba/axi4/Xbar.scala:272:23
      xbar_readys_mask_7 <= 4'hF;	// src/main/scala/tilelink/Arbiter.scala:23:23
      xbar_state_7_0 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_7_1 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_7_2 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
      xbar_state_7_3 <= 1'h0;	// src/main/scala/amba/axi4/Xbar.scala:291:24
    end
    else begin
      automatic logic xbar_ = xbar_out_0_aw_ready & xbar_out_0_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, src/main/scala/chisel3/util/Decoupled.scala:52:35
      automatic logic xbar__0 = xbar_out_1_aw_ready & xbar_out_1_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, src/main/scala/chisel3/util/Decoupled.scala:52:35
      automatic logic xbar__1 = xbar_out_2_aw_ready & xbar_out_2_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, src/main/scala/chisel3/util/Decoupled.scala:52:35
      automatic logic xbar__2 = xbar_out_3_aw_ready & xbar_out_3_aw_valid;	// src/main/scala/amba/axi4/Xbar.scala:178:19, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_awIn_0_do_enq)	// src/main/scala/chisel3/util/Decoupled.scala:264:27
        xbar_awIn_0_enq_ptr_value <= xbar_awIn_0_enq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (xbar_awIn_0_do_deq)	// src/main/scala/chisel3/util/Decoupled.scala:265:27
        xbar_awIn_0_deq_ptr_value <= xbar_awIn_0_deq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (~(xbar_awIn_0_do_enq == xbar_awIn_0_do_deq))	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27, :265:27, :277:{15,27}, :278:16
        xbar_awIn_0_maybe_full <= xbar_awIn_0_do_enq;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27
      if (xbar_awIn_1_do_enq)	// src/main/scala/chisel3/util/Decoupled.scala:264:27
        xbar_awIn_1_enq_ptr_value <= xbar_awIn_1_enq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (xbar_awIn_1_do_deq)	// src/main/scala/chisel3/util/Decoupled.scala:265:27
        xbar_awIn_1_deq_ptr_value <= xbar_awIn_1_deq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (~(xbar_awIn_1_do_enq == xbar_awIn_1_do_deq))	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27, :265:27, :277:{15,27}, :278:16
        xbar_awIn_1_maybe_full <= xbar_awIn_1_do_enq;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27
      if (xbar_awOut_0_do_enq)	// src/main/scala/chisel3/util/Decoupled.scala:264:27
        xbar_awOut_0_enq_ptr_value <= xbar_awOut_0_enq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (xbar_awOut_0_do_deq)	// src/main/scala/chisel3/util/Decoupled.scala:265:27
        xbar_awOut_0_deq_ptr_value <= xbar_awOut_0_deq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (~(xbar_awOut_0_do_enq == xbar_awOut_0_do_deq))	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27, :265:27, :277:{15,27}, :278:16
        xbar_awOut_0_maybe_full <= xbar_awOut_0_do_enq;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27
      if (xbar_awOut_1_do_enq)	// src/main/scala/chisel3/util/Decoupled.scala:264:27
        xbar_awOut_1_enq_ptr_value <= xbar_awOut_1_enq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (xbar_awOut_1_do_deq)	// src/main/scala/chisel3/util/Decoupled.scala:265:27
        xbar_awOut_1_deq_ptr_value <= xbar_awOut_1_deq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (~(xbar_awOut_1_do_enq == xbar_awOut_1_do_deq))	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27, :265:27, :277:{15,27}, :278:16
        xbar_awOut_1_maybe_full <= xbar_awOut_1_do_enq;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27
      if (xbar_awOut_2_do_enq)	// src/main/scala/chisel3/util/Decoupled.scala:264:27
        xbar_awOut_2_enq_ptr_value <= xbar_awOut_2_enq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (xbar_awOut_2_do_deq)	// src/main/scala/chisel3/util/Decoupled.scala:265:27
        xbar_awOut_2_deq_ptr_value <= xbar_awOut_2_deq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (~(xbar_awOut_2_do_enq == xbar_awOut_2_do_deq))	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27, :265:27, :277:{15,27}, :278:16
        xbar_awOut_2_maybe_full <= xbar_awOut_2_do_enq;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27
      if (xbar_awOut_3_do_enq)	// src/main/scala/chisel3/util/Decoupled.scala:264:27
        xbar_awOut_3_enq_ptr_value <= xbar_awOut_3_enq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (xbar_awOut_3_do_deq)	// src/main/scala/chisel3/util/Decoupled.scala:265:27
        xbar_awOut_3_deq_ptr_value <= xbar_awOut_3_deq_ptr_value - 1'h1;	// src/main/scala/chisel3/util/Counter.scala:61:40, :77:24
      if (~(xbar_awOut_3_do_enq == xbar_awOut_3_do_deq))	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27, :265:27, :277:{15,27}, :278:16
        xbar_awOut_3_maybe_full <= xbar_awOut_3_do_enq;	// src/main/scala/chisel3/util/Decoupled.scala:260:27, :264:27
      xbar_arFIFOMap_0_count <=
        xbar_arFIFOMap_0_count + {2'h0, xbar__arFIFOMap_0_T}
        - {2'h0, xbar__arFIFOMap_0_T_4};	// src/main/scala/amba/axi4/Xbar.scala:128:34, :130:{30,48}, :144:43, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_awFIFOMap_0_count <=
        xbar_awFIFOMap_0_count + {2'h0, xbar__awFIFOMap_0_T}
        - {2'h0, xbar__awFIFOMap_0_T_2};	// src/main/scala/amba/axi4/Xbar.scala:128:34, :130:{30,48}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_latched <=
        ~(xbar_in_0_aw_ready & xbar_in_0_aw_valid)
        & (xbar_awIn_0_io_enq_ready & xbar_awIn_0_io_enq_valid | xbar_latched);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :161:30, :165:{36,46}, :166:{30,40}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_arFIFOMap_2_count <=
        xbar_arFIFOMap_2_count + {2'h0, xbar__arFIFOMap_2_T_2}
        - {2'h0, xbar__arFIFOMap_2_T_6};	// src/main/scala/amba/axi4/Xbar.scala:128:34, :130:{30,48}, :143:25, :144:{24,43}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_awFIFOMap_2_count <=
        xbar_awFIFOMap_2_count + {2'h0, xbar__awFIFOMap_2_T_2}
        - {2'h0, xbar__awFIFOMap_2_T_5};	// src/main/scala/amba/axi4/Xbar.scala:128:34, :130:{30,48}, :147:25, :148:24, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_latched_1 <=
        ~(xbar_in_1_aw_ready & xbar_in_1_aw_valid)
        & (xbar_awIn_1_io_enq_ready & xbar_awIn_1_io_enq_valid | xbar_latched_1);	// src/main/scala/amba/axi4/Xbar.scala:90:18, :161:30, :165:{36,46}, :166:{30,40}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_latched_2 <=
        ~xbar_ & (xbar_awOut_0_io_enq_ready & xbar_awOut_0_io_enq_valid | xbar_latched_2);	// src/main/scala/amba/axi4/Xbar.scala:186:30, :190:{37,47}, :191:{31,41}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_latched_3 <=
        ~xbar__0
        & (xbar_awOut_1_io_enq_ready & xbar_awOut_1_io_enq_valid | xbar_latched_3);	// src/main/scala/amba/axi4/Xbar.scala:186:30, :190:{37,47}, :191:{31,41}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_latched_4 <=
        ~xbar__1
        & (xbar_awOut_2_io_enq_ready & xbar_awOut_2_io_enq_valid | xbar_latched_4);	// src/main/scala/amba/axi4/Xbar.scala:186:30, :190:{37,47}, :191:{31,41}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_latched_5 <=
        ~xbar__2
        & (xbar_awOut_3_io_enq_ready & xbar_awOut_3_io_enq_valid | xbar_latched_5);	// src/main/scala/amba/axi4/Xbar.scala:186:30, :190:{37,47}, :191:{31,41}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_awOut_0_io_enq_bits_idle <=
        xbar_ | ~xbar_awOut_0_io_enq_bits_anyValid & xbar_awOut_0_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_awOut_0_io_enq_bits_idle & (|xbar_awOut_0_io_enq_bits_readys_valid)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__awOut_0_io_enq_bits_readys_mask_T =
          xbar_awOut_0_io_enq_bits_readys_readys & xbar_awOut_0_io_enq_bits_readys_valid;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_awOut_0_io_enq_bits_readys_mask <=
          xbar__awOut_0_io_enq_bits_readys_mask_T
          | {xbar__awOut_0_io_enq_bits_readys_mask_T[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_awOut_0_io_enq_bits_state_0 <= xbar_awOut_0_io_enq_bits_muxState_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_awOut_0_io_enq_bits_state_1 <= xbar_awOut_0_io_enq_bits_muxState_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle <= xbar_out_0_ar_ready & xbar_out_0_ar_valid | ~xbar_anyValid & xbar_idle;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle & (|xbar_readys_valid)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__readys_mask_T =
          xbar_readys_readys & xbar_readys_valid;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_readys_mask <= xbar__readys_mask_T | {xbar__readys_mask_T[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_0 <= xbar_muxState_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_1 <= xbar_muxState_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_awOut_1_io_enq_bits_idle <=
        xbar__0 | ~xbar_awOut_1_io_enq_bits_anyValid & xbar_awOut_1_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_awOut_1_io_enq_bits_idle & (|xbar_awOut_1_io_enq_bits_readys_valid)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__awOut_1_io_enq_bits_readys_mask_T =
          xbar_awOut_1_io_enq_bits_readys_readys & xbar_awOut_1_io_enq_bits_readys_valid;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_awOut_1_io_enq_bits_readys_mask <=
          xbar__awOut_1_io_enq_bits_readys_mask_T
          | {xbar__awOut_1_io_enq_bits_readys_mask_T[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_awOut_1_io_enq_bits_state_0 <= xbar_awOut_1_io_enq_bits_muxState_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_awOut_1_io_enq_bits_state_1 <= xbar_awOut_1_io_enq_bits_muxState_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle_1 <=
        xbar_out_1_ar_ready & xbar_out_1_ar_valid | ~xbar_anyValid_1 & xbar_idle_1;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle_1 & (|xbar_readys_valid_1)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__readys_mask_T_5 =
          xbar_readys_readys_1 & xbar_readys_valid_1;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_readys_mask_1 <= xbar__readys_mask_T_5 | {xbar__readys_mask_T_5[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_1_0 <= xbar_muxState_1_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_1_1 <= xbar_muxState_1_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_awOut_2_io_enq_bits_idle <=
        xbar__1 | ~xbar_awOut_2_io_enq_bits_anyValid & xbar_awOut_2_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_awOut_2_io_enq_bits_idle & (|xbar_awOut_2_io_enq_bits_readys_valid)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__awOut_2_io_enq_bits_readys_mask_T =
          xbar_awOut_2_io_enq_bits_readys_readys & xbar_awOut_2_io_enq_bits_readys_valid;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_awOut_2_io_enq_bits_readys_mask <=
          xbar__awOut_2_io_enq_bits_readys_mask_T
          | {xbar__awOut_2_io_enq_bits_readys_mask_T[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_awOut_2_io_enq_bits_state_0 <= xbar_awOut_2_io_enq_bits_muxState_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_awOut_2_io_enq_bits_state_1 <= xbar_awOut_2_io_enq_bits_muxState_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle_2 <=
        xbar_out_2_ar_ready & xbar_out_2_ar_valid | ~xbar_anyValid_2 & xbar_idle_2;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle_2 & (|xbar_readys_valid_2)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__readys_mask_T_10 =
          xbar_readys_readys_2 & xbar_readys_valid_2;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_readys_mask_2 <= xbar__readys_mask_T_10 | {xbar__readys_mask_T_10[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_2_0 <= xbar_muxState_2_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_2_1 <= xbar_muxState_2_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_awOut_3_io_enq_bits_idle <=
        xbar__2 | ~xbar_awOut_3_io_enq_bits_anyValid & xbar_awOut_3_io_enq_bits_idle;	// src/main/scala/amba/axi4/Xbar.scala:272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_awOut_3_io_enq_bits_idle & (|xbar_awOut_3_io_enq_bits_readys_valid)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__awOut_3_io_enq_bits_readys_mask_T =
          xbar_awOut_3_io_enq_bits_readys_readys & xbar_awOut_3_io_enq_bits_readys_valid;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_awOut_3_io_enq_bits_readys_mask <=
          xbar__awOut_3_io_enq_bits_readys_mask_T
          | {xbar__awOut_3_io_enq_bits_readys_mask_T[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_awOut_3_io_enq_bits_state_0 <= xbar_awOut_3_io_enq_bits_muxState_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_awOut_3_io_enq_bits_state_1 <= xbar_awOut_3_io_enq_bits_muxState_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle_3 <=
        xbar_out_3_ar_ready & xbar_out_3_ar_valid | ~xbar_anyValid_3 & xbar_idle_3;	// src/main/scala/amba/axi4/Xbar.scala:178:19, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle_3 & (|xbar_readys_valid_3)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [1:0] xbar__readys_mask_T_15 =
          xbar_readys_readys_3 & xbar_readys_valid_3;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        xbar_readys_mask_3 <= xbar__readys_mask_T_15 | {xbar__readys_mask_T_15[0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, :28:29, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_3_0 <= xbar_muxState_3_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_3_1 <= xbar_muxState_3_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle_4 <=
        xbar_in_0_r_ready & xbar_in_0_r_valid | ~xbar_anyValid_4 & xbar_idle_4;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle_4 & (|xbar_readys_valid_4)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [3:0] xbar__readys_mask_T_20 =
          xbar_readys_readys_4 & xbar_readys_valid_4;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        automatic logic [3:0] xbar__readys_mask_T_23 =
          xbar__readys_mask_T_20 | {xbar__readys_mask_T_20[2:0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:28:29, src/main/scala/util/package.scala:253:{43,53}
        xbar_readys_mask_4 <=
          xbar__readys_mask_T_23 | {xbar__readys_mask_T_23[1:0], 2'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_4_0 <= xbar_muxState_4_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_4_1 <= xbar_muxState_4_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_4_2 <= xbar_muxState_4_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_4_3 <= xbar_muxState_4_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle_5 <=
        xbar_in_0_b_ready & xbar_in_0_b_valid | ~xbar_anyValid_5 & xbar_idle_5;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle_5 & (|xbar_readys_valid_5)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [3:0] xbar__readys_mask_T_28 =
          xbar_readys_readys_5 & xbar_readys_valid_5;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        automatic logic [3:0] xbar__readys_mask_T_31 =
          xbar__readys_mask_T_28 | {xbar__readys_mask_T_28[2:0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:28:29, src/main/scala/util/package.scala:253:{43,53}
        xbar_readys_mask_5 <=
          xbar__readys_mask_T_31 | {xbar__readys_mask_T_31[1:0], 2'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_5_0 <= xbar_muxState_5_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_5_1 <= xbar_muxState_5_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_5_2 <= xbar_muxState_5_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_5_3 <= xbar_muxState_5_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle_6 <=
        xbar_in_1_r_ready & xbar_in_1_r_valid | ~xbar_anyValid_6 & xbar_idle_6;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle_6 & (|xbar_readys_valid_6)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [3:0] xbar__readys_mask_T_36 =
          xbar_readys_readys_6 & xbar_readys_valid_6;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        automatic logic [3:0] xbar__readys_mask_T_39 =
          xbar__readys_mask_T_36 | {xbar__readys_mask_T_36[2:0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:28:29, src/main/scala/util/package.scala:253:{43,53}
        xbar_readys_mask_6 <=
          xbar__readys_mask_T_39 | {xbar__readys_mask_T_39[1:0], 2'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_6_0 <= xbar_muxState_6_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_6_1 <= xbar_muxState_6_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_6_2 <= xbar_muxState_6_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_6_3 <= xbar_muxState_6_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_idle_7 <=
        xbar_in_1_b_ready & xbar_in_1_b_valid | ~xbar_anyValid_7 & xbar_idle_7;	// src/main/scala/amba/axi4/Xbar.scala:90:18, :272:23, :276:36, :296:{21,28}, :297:{22,29}, src/main/scala/chisel3/util/Decoupled.scala:52:35
      if (xbar_idle_7 & (|xbar_readys_valid_7)) begin	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:21:23, :27:{18,27}
        automatic logic [3:0] xbar__readys_mask_T_44 =
          xbar_readys_readys_7 & xbar_readys_valid_7;	// src/main/scala/tilelink/Arbiter.scala:21:23, :26:18, :28:29
        automatic logic [3:0] xbar__readys_mask_T_47 =
          xbar__readys_mask_T_44 | {xbar__readys_mask_T_44[2:0], 1'h0};	// src/main/scala/tilelink/Arbiter.scala:28:29, src/main/scala/util/package.scala:253:{43,53}
        xbar_readys_mask_7 <=
          xbar__readys_mask_T_47 | {xbar__readys_mask_T_47[1:0], 2'h0};	// src/main/scala/tilelink/Arbiter.scala:23:23, src/main/scala/util/package.scala:253:{43,53}
      end
      xbar_state_7_0 <= xbar_muxState_7_0;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_7_1 <= xbar_muxState_7_1;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_7_2 <= xbar_muxState_7_2;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
      xbar_state_7_3 <= xbar_muxState_7_3;	// src/main/scala/amba/axi4/Xbar.scala:291:24, :292:23
    end
    if (xbar__arFIFOMap_0_T)	// src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_arFIFOMap_0_last <= xbar_arTag;	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/chisel3/util/OneHot.scala:32:10
    if (xbar__awFIFOMap_0_T)	// src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_awFIFOMap_0_last <= xbar_awTag;	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/chisel3/util/OneHot.scala:32:10
    if (xbar__arFIFOMap_2_T_2)	// src/main/scala/amba/axi4/Xbar.scala:143:25, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_arFIFOMap_2_last <= xbar_arTag_1;	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/chisel3/util/OneHot.scala:32:10
    if (xbar__awFIFOMap_2_T_2)	// src/main/scala/amba/axi4/Xbar.scala:147:25, src/main/scala/chisel3/util/Decoupled.scala:52:35
      xbar_awFIFOMap_2_last <= xbar_awTag_1;	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/chisel3/util/OneHot.scala:32:10
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    initial begin
      automatic logic [31:0] _RANDOM[0:3];
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [2:0] i = 3'h0; i < 3'h4; i += 3'h1) begin
          _RANDOM[i[1:0]] = `RANDOM;
        end
        xbar_awIn_0_enq_ptr_value = _RANDOM[2'h0][0];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awIn_0_deq_ptr_value = _RANDOM[2'h0][1];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awIn_0_maybe_full = _RANDOM[2'h0][2];	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:260:27
        xbar_awIn_1_enq_ptr_value = _RANDOM[2'h0][3];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awIn_1_deq_ptr_value = _RANDOM[2'h0][4];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awIn_1_maybe_full = _RANDOM[2'h0][5];	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:260:27
        xbar_awOut_0_enq_ptr_value = _RANDOM[2'h0][6];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_0_deq_ptr_value = _RANDOM[2'h0][7];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_0_maybe_full = _RANDOM[2'h0][8];	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:260:27
        xbar_awOut_1_enq_ptr_value = _RANDOM[2'h0][9];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_1_deq_ptr_value = _RANDOM[2'h0][10];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_1_maybe_full = _RANDOM[2'h0][11];	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:260:27
        xbar_awOut_2_enq_ptr_value = _RANDOM[2'h0][12];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_2_deq_ptr_value = _RANDOM[2'h0][13];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_2_maybe_full = _RANDOM[2'h0][14];	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:260:27
        xbar_awOut_3_enq_ptr_value = _RANDOM[2'h0][15];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_3_deq_ptr_value = _RANDOM[2'h0][16];	// src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awOut_3_maybe_full = _RANDOM[2'h0][17];	// src/main/scala/chisel3/util/Counter.scala:61:40, src/main/scala/chisel3/util/Decoupled.scala:260:27
        xbar_arFIFOMap_0_count = _RANDOM[2'h0][20:18];	// src/main/scala/amba/axi4/Xbar.scala:128:34, src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_arFIFOMap_0_last = _RANDOM[2'h0][22:21];	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awFIFOMap_0_count = _RANDOM[2'h0][25:23];	// src/main/scala/amba/axi4/Xbar.scala:128:34, src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_awFIFOMap_0_last = _RANDOM[2'h0][27:26];	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_latched = _RANDOM[2'h0][28];	// src/main/scala/amba/axi4/Xbar.scala:161:30, src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_arFIFOMap_2_count = _RANDOM[2'h0][31:29];	// src/main/scala/amba/axi4/Xbar.scala:128:34, src/main/scala/chisel3/util/Counter.scala:61:40
        xbar_arFIFOMap_2_last = _RANDOM[2'h1][1:0];	// src/main/scala/amba/axi4/Xbar.scala:129:29
        xbar_awFIFOMap_2_count = _RANDOM[2'h1][4:2];	// src/main/scala/amba/axi4/Xbar.scala:128:34, :129:29
        xbar_awFIFOMap_2_last = _RANDOM[2'h1][6:5];	// src/main/scala/amba/axi4/Xbar.scala:129:29
        xbar_latched_1 = _RANDOM[2'h1][7];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :161:30
        xbar_latched_2 = _RANDOM[2'h1][8];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :186:30
        xbar_latched_3 = _RANDOM[2'h1][9];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :186:30
        xbar_latched_4 = _RANDOM[2'h1][10];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :186:30
        xbar_latched_5 = _RANDOM[2'h1][11];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :186:30
        xbar_awOut_0_io_enq_bits_idle = _RANDOM[2'h1][12];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :272:23
        xbar_awOut_0_io_enq_bits_readys_mask = _RANDOM[2'h1][14:13];	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_awOut_0_io_enq_bits_state_0 = _RANDOM[2'h1][15];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_awOut_0_io_enq_bits_state_1 = _RANDOM[2'h1][16];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_idle = _RANDOM[2'h1][17];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :272:23
        xbar_readys_mask = _RANDOM[2'h1][19:18];	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_0 = _RANDOM[2'h1][20];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_state_1 = _RANDOM[2'h1][21];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_awOut_1_io_enq_bits_idle = _RANDOM[2'h1][22];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :272:23
        xbar_awOut_1_io_enq_bits_readys_mask = _RANDOM[2'h1][24:23];	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_awOut_1_io_enq_bits_state_0 = _RANDOM[2'h1][25];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_awOut_1_io_enq_bits_state_1 = _RANDOM[2'h1][26];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_idle_1 = _RANDOM[2'h1][27];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :272:23
        xbar_readys_mask_1 = _RANDOM[2'h1][29:28];	// src/main/scala/amba/axi4/Xbar.scala:129:29, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_1_0 = _RANDOM[2'h1][30];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_state_1_1 = _RANDOM[2'h1][31];	// src/main/scala/amba/axi4/Xbar.scala:129:29, :291:24
        xbar_awOut_2_io_enq_bits_idle = _RANDOM[2'h2][0];	// src/main/scala/amba/axi4/Xbar.scala:272:23
        xbar_awOut_2_io_enq_bits_readys_mask = _RANDOM[2'h2][2:1];	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_awOut_2_io_enq_bits_state_0 = _RANDOM[2'h2][3];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_awOut_2_io_enq_bits_state_1 = _RANDOM[2'h2][4];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_idle_2 = _RANDOM[2'h2][5];	// src/main/scala/amba/axi4/Xbar.scala:272:23
        xbar_readys_mask_2 = _RANDOM[2'h2][7:6];	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_2_0 = _RANDOM[2'h2][8];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_state_2_1 = _RANDOM[2'h2][9];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_awOut_3_io_enq_bits_idle = _RANDOM[2'h2][10];	// src/main/scala/amba/axi4/Xbar.scala:272:23
        xbar_awOut_3_io_enq_bits_readys_mask = _RANDOM[2'h2][12:11];	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_awOut_3_io_enq_bits_state_0 = _RANDOM[2'h2][13];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_awOut_3_io_enq_bits_state_1 = _RANDOM[2'h2][14];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_idle_3 = _RANDOM[2'h2][15];	// src/main/scala/amba/axi4/Xbar.scala:272:23
        xbar_readys_mask_3 = _RANDOM[2'h2][17:16];	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_3_0 = _RANDOM[2'h2][18];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_state_3_1 = _RANDOM[2'h2][19];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_idle_4 = _RANDOM[2'h2][20];	// src/main/scala/amba/axi4/Xbar.scala:272:23
        xbar_readys_mask_4 = _RANDOM[2'h2][24:21];	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_4_0 = _RANDOM[2'h2][25];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_state_4_1 = _RANDOM[2'h2][26];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_state_4_2 = _RANDOM[2'h2][27];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_state_4_3 = _RANDOM[2'h2][28];	// src/main/scala/amba/axi4/Xbar.scala:272:23, :291:24
        xbar_idle_5 = _RANDOM[2'h2][29];	// src/main/scala/amba/axi4/Xbar.scala:272:23
        xbar_readys_mask_5 = {_RANDOM[2'h2][31:30], _RANDOM[2'h3][1:0]};	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_5_0 = _RANDOM[2'h3][2];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_5_1 = _RANDOM[2'h3][3];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_5_2 = _RANDOM[2'h3][4];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_5_3 = _RANDOM[2'h3][5];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_idle_6 = _RANDOM[2'h3][6];	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_readys_mask_6 = _RANDOM[2'h3][10:7];	// src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_6_0 = _RANDOM[2'h3][11];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_6_1 = _RANDOM[2'h3][12];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_6_2 = _RANDOM[2'h3][13];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_6_3 = _RANDOM[2'h3][14];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_idle_7 = _RANDOM[2'h3][15];	// src/main/scala/amba/axi4/Xbar.scala:272:23, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_readys_mask_7 = _RANDOM[2'h3][19:16];	// src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_7_0 = _RANDOM[2'h3][20];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_7_1 = _RANDOM[2'h3][21];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_7_2 = _RANDOM[2'h3][22];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
        xbar_state_7_3 = _RANDOM[2'h3][23];	// src/main/scala/amba/axi4/Xbar.scala:291:24, src/main/scala/tilelink/Arbiter.scala:23:23
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  ram_2x4 ram_ext (	// src/main/scala/chisel3/util/Decoupled.scala:257:91
    .R0_addr (xbar_awIn_0_deq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R0_data (_ram_ext_R0_data_4),
    .W0_addr (xbar_awIn_0_enq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .W0_en   (xbar_awIn_0_do_enq),	// src/main/scala/chisel3/util/Decoupled.scala:264:27
    .W0_clk  (clock),
    .W0_data (xbar_awIn_0_io_enq_bits)
  );	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  ram_2x4 ram_ext_0 (	// src/main/scala/chisel3/util/Decoupled.scala:257:91
    .R0_addr (xbar_awIn_1_deq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R0_data (_ram_ext_R0_data_3),
    .W0_addr (xbar_awIn_1_enq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .W0_en   (xbar_awIn_1_do_enq),	// src/main/scala/chisel3/util/Decoupled.scala:264:27
    .W0_clk  (clock),
    .W0_data (xbar_awIn_1_io_enq_bits)
  );	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  ram_2x2 ram_ext_1 (	// src/main/scala/chisel3/util/Decoupled.scala:257:91
    .R0_addr (xbar_awOut_0_deq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R0_data (_ram_ext_R0_data_2),
    .W0_addr (xbar_awOut_0_enq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .W0_en   (xbar_awOut_0_do_enq),	// src/main/scala/chisel3/util/Decoupled.scala:264:27
    .W0_clk  (clock),
    .W0_data (xbar_awOut_0_io_enq_bits)
  );	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  ram_2x2 ram_ext_2 (	// src/main/scala/chisel3/util/Decoupled.scala:257:91
    .R0_addr (xbar_awOut_1_deq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R0_data (_ram_ext_R0_data_1),
    .W0_addr (xbar_awOut_1_enq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .W0_en   (xbar_awOut_1_do_enq),	// src/main/scala/chisel3/util/Decoupled.scala:264:27
    .W0_clk  (clock),
    .W0_data (xbar_awOut_1_io_enq_bits)
  );	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  ram_2x2 ram_ext_3 (	// src/main/scala/chisel3/util/Decoupled.scala:257:91
    .R0_addr (xbar_awOut_2_deq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R0_data (_ram_ext_R0_data_0),
    .W0_addr (xbar_awOut_2_enq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .W0_en   (xbar_awOut_2_do_enq),	// src/main/scala/chisel3/util/Decoupled.scala:264:27
    .W0_clk  (clock),
    .W0_data (xbar_awOut_2_io_enq_bits)
  );	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  ram_2x2 ram_ext_4 (	// src/main/scala/chisel3/util/Decoupled.scala:257:91
    .R0_addr (xbar_awOut_3_deq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .R0_en   (1'h1),
    .R0_clk  (clock),
    .R0_data (_ram_ext_R0_data),
    .W0_addr (xbar_awOut_3_enq_ptr_value),	// src/main/scala/chisel3/util/Counter.scala:61:40
    .W0_en   (xbar_awOut_3_do_enq),	// src/main/scala/chisel3/util/Decoupled.scala:264:27
    .W0_clk  (clock),
    .W0_data (xbar_awOut_3_io_enq_bits)
  );	// src/main/scala/chisel3/util/Decoupled.scala:257:91
  assign master1_aw_ready = master1_aw_ready_0;
  assign master1_w_ready = master1_w_ready_0;
  assign master1_b_valid = master1_b_valid_0;
  assign master1_b_bits_id = 8'h0;
  assign master1_b_bits_resp = master1_b_bits_resp_0;
  assign master1_ar_ready = master1_ar_ready_0;
  assign master1_r_valid = master1_r_valid_0;
  assign master1_r_bits_id = 8'h0;
  assign master1_r_bits_data = master1_r_bits_data_0;
  assign master1_r_bits_resp = master1_r_bits_resp_0;
  assign master1_r_bits_last = master1_r_bits_last_0;
  assign master2_aw_ready = master2_aw_ready_0;
  assign master2_w_ready = master2_w_ready_0;
  assign master2_b_valid = master2_b_valid_0;
  assign master2_b_bits_id = master2_b_bits_id_0;
  assign master2_b_bits_resp = master2_b_bits_resp_0;
  assign master2_ar_ready = master2_ar_ready_0;
  assign master2_r_valid = master2_r_valid_0;
  assign master2_r_bits_id = master2_r_bits_id_0;
  assign master2_r_bits_data = master2_r_bits_data_0;
  assign master2_r_bits_resp = master2_r_bits_resp_0;
  assign master2_r_bits_last = master2_r_bits_last_0;
  assign slave1_aw_valid = slave1_aw_valid_0;
  assign slave1_aw_bits_id = slave1_aw_bits_id_0;
  assign slave1_aw_bits_addr = slave1_aw_bits_addr_0;
  assign slave1_aw_bits_len = slave1_aw_bits_len_0;
  assign slave1_aw_bits_size = slave1_aw_bits_size_0;
  assign slave1_aw_bits_burst = slave1_aw_bits_burst_0;
  assign slave1_aw_bits_lock = slave1_aw_bits_lock_0;
  assign slave1_aw_bits_cache = slave1_aw_bits_cache_0;
  assign slave1_aw_bits_prot = slave1_aw_bits_prot_0;
  assign slave1_aw_bits_qos = slave1_aw_bits_qos_0;
  assign slave1_w_valid = slave1_w_valid_0;
  assign slave1_w_bits_data = slave1_w_bits_data_0;
  assign slave1_w_bits_strb = slave1_w_bits_strb_0;
  assign slave1_w_bits_last = slave1_w_bits_last_0;
  assign slave1_b_ready = slave1_b_ready_0;
  assign slave1_ar_valid = slave1_ar_valid_0;
  assign slave1_ar_bits_id = slave1_ar_bits_id_0;
  assign slave1_ar_bits_addr = slave1_ar_bits_addr_0;
  assign slave1_ar_bits_len = slave1_ar_bits_len_0;
  assign slave1_ar_bits_size = slave1_ar_bits_size_0;
  assign slave1_ar_bits_burst = slave1_ar_bits_burst_0;
  assign slave1_ar_bits_lock = slave1_ar_bits_lock_0;
  assign slave1_ar_bits_cache = slave1_ar_bits_cache_0;
  assign slave1_ar_bits_prot = slave1_ar_bits_prot_0;
  assign slave1_ar_bits_qos = slave1_ar_bits_qos_0;
  assign slave1_r_ready = slave1_r_ready_0;
  assign slave2_aw_valid = slave2_aw_valid_0;
  assign slave2_aw_bits_id = slave2_aw_bits_id_0;
  assign slave2_aw_bits_addr = slave2_aw_bits_addr_0;
  assign slave2_aw_bits_len = slave2_aw_bits_len_0;
  assign slave2_aw_bits_size = slave2_aw_bits_size_0;
  assign slave2_aw_bits_burst = slave2_aw_bits_burst_0;
  assign slave2_aw_bits_lock = slave2_aw_bits_lock_0;
  assign slave2_aw_bits_cache = slave2_aw_bits_cache_0;
  assign slave2_aw_bits_prot = slave2_aw_bits_prot_0;
  assign slave2_aw_bits_qos = slave2_aw_bits_qos_0;
  assign slave2_w_valid = slave2_w_valid_0;
  assign slave2_w_bits_data = slave2_w_bits_data_0;
  assign slave2_w_bits_strb = slave2_w_bits_strb_0;
  assign slave2_w_bits_last = slave2_w_bits_last_0;
  assign slave2_b_ready = slave2_b_ready_0;
  assign slave2_ar_valid = slave2_ar_valid_0;
  assign slave2_ar_bits_id = slave2_ar_bits_id_0;
  assign slave2_ar_bits_addr = slave2_ar_bits_addr_0;
  assign slave2_ar_bits_len = slave2_ar_bits_len_0;
  assign slave2_ar_bits_size = slave2_ar_bits_size_0;
  assign slave2_ar_bits_burst = slave2_ar_bits_burst_0;
  assign slave2_ar_bits_lock = slave2_ar_bits_lock_0;
  assign slave2_ar_bits_cache = slave2_ar_bits_cache_0;
  assign slave2_ar_bits_prot = slave2_ar_bits_prot_0;
  assign slave2_ar_bits_qos = slave2_ar_bits_qos_0;
  assign slave2_r_ready = slave2_r_ready_0;
  assign slave3_aw_valid = slave3_aw_valid_0;
  assign slave3_aw_bits_id = slave3_aw_bits_id_0;
  assign slave3_aw_bits_addr = slave3_aw_bits_addr_0;
  assign slave3_aw_bits_len = slave3_aw_bits_len_0;
  assign slave3_aw_bits_size = slave3_aw_bits_size_0;
  assign slave3_aw_bits_burst = slave3_aw_bits_burst_0;
  assign slave3_aw_bits_lock = slave3_aw_bits_lock_0;
  assign slave3_aw_bits_cache = slave3_aw_bits_cache_0;
  assign slave3_aw_bits_prot = slave3_aw_bits_prot_0;
  assign slave3_aw_bits_qos = slave3_aw_bits_qos_0;
  assign slave3_w_valid = slave3_w_valid_0;
  assign slave3_w_bits_data = slave3_w_bits_data_0;
  assign slave3_w_bits_strb = slave3_w_bits_strb_0;
  assign slave3_w_bits_last = slave3_w_bits_last_0;
  assign slave3_b_ready = slave3_b_ready_0;
  assign slave3_ar_valid = slave3_ar_valid_0;
  assign slave3_ar_bits_id = slave3_ar_bits_id_0;
  assign slave3_ar_bits_addr = slave3_ar_bits_addr_0;
  assign slave3_ar_bits_len = slave3_ar_bits_len_0;
  assign slave3_ar_bits_size = slave3_ar_bits_size_0;
  assign slave3_ar_bits_burst = slave3_ar_bits_burst_0;
  assign slave3_ar_bits_lock = slave3_ar_bits_lock_0;
  assign slave3_ar_bits_cache = slave3_ar_bits_cache_0;
  assign slave3_ar_bits_prot = slave3_ar_bits_prot_0;
  assign slave3_ar_bits_qos = slave3_ar_bits_qos_0;
  assign slave3_r_ready = slave3_r_ready_0;
  assign slave4_aw_valid = slave4_aw_valid_0;
  assign slave4_aw_bits_id = slave4_aw_bits_id_0;
  assign slave4_aw_bits_addr = slave4_aw_bits_addr_0;
  assign slave4_aw_bits_len = slave4_aw_bits_len_0;
  assign slave4_aw_bits_size = slave4_aw_bits_size_0;
  assign slave4_aw_bits_burst = slave4_aw_bits_burst_0;
  assign slave4_aw_bits_lock = slave4_aw_bits_lock_0;
  assign slave4_aw_bits_cache = slave4_aw_bits_cache_0;
  assign slave4_aw_bits_prot = slave4_aw_bits_prot_0;
  assign slave4_aw_bits_qos = slave4_aw_bits_qos_0;
  assign slave4_w_valid = slave4_w_valid_0;
  assign slave4_w_bits_data = slave4_w_bits_data_0;
  assign slave4_w_bits_strb = slave4_w_bits_strb_0;
  assign slave4_w_bits_last = slave4_w_bits_last_0;
  assign slave4_b_ready = slave4_b_ready_0;
  assign slave4_ar_valid = slave4_ar_valid_0;
  assign slave4_ar_bits_id = slave4_ar_bits_id_0;
  assign slave4_ar_bits_addr = slave4_ar_bits_addr_0;
  assign slave4_ar_bits_len = slave4_ar_bits_len_0;
  assign slave4_ar_bits_size = slave4_ar_bits_size_0;
  assign slave4_ar_bits_burst = slave4_ar_bits_burst_0;
  assign slave4_ar_bits_lock = slave4_ar_bits_lock_0;
  assign slave4_ar_bits_cache = slave4_ar_bits_cache_0;
  assign slave4_ar_bits_prot = slave4_ar_bits_prot_0;
  assign slave4_ar_bits_qos = slave4_ar_bits_qos_0;
  assign slave4_r_ready = slave4_r_ready_0;
endmodule


        
/* verilator lint_off WIDTH */        
module AXI4XBar2x4 
   (
   input logic  clock,
   input logic  reset,
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION.inward master1,
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION.inward master2,
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION.outward slave1,
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION.outward slave2,
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION.outward slave3,
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION.outward slave4
   );

   


    AXI4XBar2x4_inner inner
      (
        .clock(clock),
        .reset(reset),
        .master1_aw_bits_id(master1.AWID),
        .master1_aw_bits_addr(master1.AWADDR),
        .master1_aw_bits_len(master1.AWLEN),
        .master1_aw_bits_size(master1.AWSIZE),
        .master1_aw_bits_burst(master1.AWBURST),
        .master1_aw_bits_lock(master1.AWLOCK),
        .master1_aw_bits_cache(master1.AWCACHE),
        .master1_aw_bits_prot(master1.AWPROT),
        .master1_aw_valid(master1.AWVALID),
        .master1_aw_ready(master1.AWREADY),
        .master1_w_bits_data(master1.WDATA),
        .master1_w_bits_strb(master1.WSTRB),
        .master1_w_bits_last(master1.WLAST),
        .master1_w_valid(master1.WVALID),
        .master1_w_ready(master1.WREADY),
        .master1_b_bits_id(master1.BID),
        .master1_b_bits_resp(master1.BRESP),
        .master1_b_valid(master1.BVALID),
        .master1_b_ready(master1.BREADY),
        .master1_ar_bits_id(master1.ARID),
        .master1_ar_bits_addr(master1.ARADDR),
        .master1_ar_bits_len(master1.ARLEN),
        .master1_ar_bits_size(master1.ARSIZE),
        .master1_ar_bits_burst(master1.ARBURST),
        .master1_ar_bits_lock(master1.ARLOCK),
        .master1_ar_bits_cache(master1.ARCACHE),
        .master1_ar_bits_prot(master1.ARPROT),
        .master1_ar_valid(master1.ARVALID),
        .master1_ar_ready(master1.ARREADY),
        .master1_r_bits_id(master1.RID),
        .master1_r_bits_data(master1.RDATA),
        .master1_r_bits_resp(master1.RRESP),
        .master1_r_bits_last(master1.RLAST),
        .master1_r_valid(master1.RVALID),
        .master1_r_ready(master1.RREADY),
        .master1_ar_bits_qos(master1.ARQOS),
        .master1_aw_bits_qos(master1.AWQOS),
        .master2_aw_bits_id(master2.AWID),
        .master2_aw_bits_addr(master2.AWADDR),
        .master2_aw_bits_len(master2.AWLEN),
        .master2_aw_bits_size(master2.AWSIZE),
        .master2_aw_bits_burst(master2.AWBURST),
        .master2_aw_bits_lock(master2.AWLOCK),
        .master2_aw_bits_cache(master2.AWCACHE),
        .master2_aw_bits_prot(master2.AWPROT),
        .master2_aw_valid(master2.AWVALID),
        .master2_aw_ready(master2.AWREADY),
        .master2_w_bits_data(master2.WDATA),
        .master2_w_bits_strb(master2.WSTRB),
        .master2_w_bits_last(master2.WLAST),
        .master2_w_valid(master2.WVALID),
        .master2_w_ready(master2.WREADY),
        .master2_b_bits_id(master2.BID),
        .master2_b_bits_resp(master2.BRESP),
        .master2_b_valid(master2.BVALID),
        .master2_b_ready(master2.BREADY),
        .master2_ar_bits_id(master2.ARID),
        .master2_ar_bits_addr(master2.ARADDR),
        .master2_ar_bits_len(master2.ARLEN),
        .master2_ar_bits_size(master2.ARSIZE),
        .master2_ar_bits_burst(master2.ARBURST),
        .master2_ar_bits_lock(master2.ARLOCK),
        .master2_ar_bits_cache(master2.ARCACHE),
        .master2_ar_bits_prot(master2.ARPROT),
        .master2_ar_valid(master2.ARVALID),
        .master2_ar_ready(master2.ARREADY),
        .master2_r_bits_id(master2.RID),
        .master2_r_bits_data(master2.RDATA),
        .master2_r_bits_resp(master2.RRESP),
        .master2_r_bits_last(master2.RLAST),
        .master2_r_valid(master2.RVALID),
        .master2_r_ready(master2.RREADY),
        .master2_ar_bits_qos(master2.ARQOS),
        .master2_aw_bits_qos(master2.AWQOS),
        .slave1_aw_bits_id(slave1.AWID),
        .slave1_aw_bits_addr(slave1.AWADDR),
        .slave1_aw_bits_len(slave1.AWLEN),
        .slave1_aw_bits_size(slave1.AWSIZE),
        .slave1_aw_bits_burst(slave1.AWBURST),
        .slave1_aw_bits_lock(slave1.AWLOCK),
        .slave1_aw_bits_cache(slave1.AWCACHE),
        .slave1_aw_bits_prot(slave1.AWPROT),
        .slave1_aw_valid(slave1.AWVALID),
        .slave1_aw_ready(slave1.AWREADY),
        .slave1_w_bits_data(slave1.WDATA),
        .slave1_w_bits_strb(slave1.WSTRB),
        .slave1_w_bits_last(slave1.WLAST),
        .slave1_w_valid(slave1.WVALID),
        .slave1_w_ready(slave1.WREADY),
        .slave1_b_bits_id(slave1.BID),
        .slave1_b_bits_resp(slave1.BRESP),
        .slave1_b_valid(slave1.BVALID),
        .slave1_b_ready(slave1.BREADY),
        .slave1_ar_bits_id(slave1.ARID),
        .slave1_ar_bits_addr(slave1.ARADDR),
        .slave1_ar_bits_len(slave1.ARLEN),
        .slave1_ar_bits_size(slave1.ARSIZE),
        .slave1_ar_bits_burst(slave1.ARBURST),
        .slave1_ar_bits_lock(slave1.ARLOCK),
        .slave1_ar_bits_cache(slave1.ARCACHE),
        .slave1_ar_bits_prot(slave1.ARPROT),
        .slave1_ar_valid(slave1.ARVALID),
        .slave1_ar_ready(slave1.ARREADY),
        .slave1_r_bits_id(slave1.RID),
        .slave1_r_bits_data(slave1.RDATA),
        .slave1_r_bits_resp(slave1.RRESP),
        .slave1_r_bits_last(slave1.RLAST),
        .slave1_r_valid(slave1.RVALID),
        .slave1_r_ready(slave1.RREADY),
        .slave1_ar_bits_qos(slave1.ARQOS),
        .slave1_aw_bits_qos(slave1.AWQOS),
        .slave2_aw_bits_id(slave2.AWID),
        .slave2_aw_bits_addr(slave2.AWADDR),
        .slave2_aw_bits_len(slave2.AWLEN),
        .slave2_aw_bits_size(slave2.AWSIZE),
        .slave2_aw_bits_burst(slave2.AWBURST),
        .slave2_aw_bits_lock(slave2.AWLOCK),
        .slave2_aw_bits_cache(slave2.AWCACHE),
        .slave2_aw_bits_prot(slave2.AWPROT),
        .slave2_aw_valid(slave2.AWVALID),
        .slave2_aw_ready(slave2.AWREADY),
        .slave2_w_bits_data(slave2.WDATA),
        .slave2_w_bits_strb(slave2.WSTRB),
        .slave2_w_bits_last(slave2.WLAST),
        .slave2_w_valid(slave2.WVALID),
        .slave2_w_ready(slave2.WREADY),
        .slave2_b_bits_id(slave2.BID),
        .slave2_b_bits_resp(slave2.BRESP),
        .slave2_b_valid(slave2.BVALID),
        .slave2_b_ready(slave2.BREADY),
        .slave2_ar_bits_id(slave2.ARID),
        .slave2_ar_bits_addr(slave2.ARADDR),
        .slave2_ar_bits_len(slave2.ARLEN),
        .slave2_ar_bits_size(slave2.ARSIZE),
        .slave2_ar_bits_burst(slave2.ARBURST),
        .slave2_ar_bits_lock(slave2.ARLOCK),
        .slave2_ar_bits_cache(slave2.ARCACHE),
        .slave2_ar_bits_prot(slave2.ARPROT),
        .slave2_ar_valid(slave2.ARVALID),
        .slave2_ar_ready(slave2.ARREADY),
        .slave2_r_bits_id(slave2.RID),
        .slave2_r_bits_data(slave2.RDATA),
        .slave2_r_bits_resp(slave2.RRESP),
        .slave2_r_bits_last(slave2.RLAST),
        .slave2_r_valid(slave2.RVALID),
        .slave2_r_ready(slave2.RREADY),
        .slave2_ar_bits_qos(slave2.ARQOS),
        .slave2_aw_bits_qos(slave2.AWQOS),
        .slave3_aw_bits_id(slave3.AWID),
        .slave3_aw_bits_addr(slave3.AWADDR),
        .slave3_aw_bits_len(slave3.AWLEN),
        .slave3_aw_bits_size(slave3.AWSIZE),
        .slave3_aw_bits_burst(slave3.AWBURST),
        .slave3_aw_bits_lock(slave3.AWLOCK),
        .slave3_aw_bits_cache(slave3.AWCACHE),
        .slave3_aw_bits_prot(slave3.AWPROT),
        .slave3_aw_valid(slave3.AWVALID),
        .slave3_aw_ready(slave3.AWREADY),
        .slave3_w_bits_data(slave3.WDATA),
        .slave3_w_bits_strb(slave3.WSTRB),
        .slave3_w_bits_last(slave3.WLAST),
        .slave3_w_valid(slave3.WVALID),
        .slave3_w_ready(slave3.WREADY),
        .slave3_b_bits_id(slave3.BID),
        .slave3_b_bits_resp(slave3.BRESP),
        .slave3_b_valid(slave3.BVALID),
        .slave3_b_ready(slave3.BREADY),
        .slave3_ar_bits_id(slave3.ARID),
        .slave3_ar_bits_addr(slave3.ARADDR),
        .slave3_ar_bits_len(slave3.ARLEN),
        .slave3_ar_bits_size(slave3.ARSIZE),
        .slave3_ar_bits_burst(slave3.ARBURST),
        .slave3_ar_bits_lock(slave3.ARLOCK),
        .slave3_ar_bits_cache(slave3.ARCACHE),
        .slave3_ar_bits_prot(slave3.ARPROT),
        .slave3_ar_valid(slave3.ARVALID),
        .slave3_ar_ready(slave3.ARREADY),
        .slave3_r_bits_id(slave3.RID),
        .slave3_r_bits_data(slave3.RDATA),
        .slave3_r_bits_resp(slave3.RRESP),
        .slave3_r_bits_last(slave3.RLAST),
        .slave3_r_valid(slave3.RVALID),
        .slave3_r_ready(slave3.RREADY),
        .slave3_ar_bits_qos(slave3.ARQOS),
        .slave3_aw_bits_qos(slave3.AWQOS),
        .slave4_aw_bits_id(slave4.AWID),
        .slave4_aw_bits_addr(slave4.AWADDR),
        .slave4_aw_bits_len(slave4.AWLEN),
        .slave4_aw_bits_size(slave4.AWSIZE),
        .slave4_aw_bits_burst(slave4.AWBURST),
        .slave4_aw_bits_lock(slave4.AWLOCK),
        .slave4_aw_bits_cache(slave4.AWCACHE),
        .slave4_aw_bits_prot(slave4.AWPROT),
        .slave4_aw_valid(slave4.AWVALID),
        .slave4_aw_ready(slave4.AWREADY),
        .slave4_w_bits_data(slave4.WDATA),
        .slave4_w_bits_strb(slave4.WSTRB),
        .slave4_w_bits_last(slave4.WLAST),
        .slave4_w_valid(slave4.WVALID),
        .slave4_w_ready(slave4.WREADY),
        .slave4_b_bits_id(slave4.BID),
        .slave4_b_bits_resp(slave4.BRESP),
        .slave4_b_valid(slave4.BVALID),
        .slave4_b_ready(slave4.BREADY),
        .slave4_ar_bits_id(slave4.ARID),
        .slave4_ar_bits_addr(slave4.ARADDR),
        .slave4_ar_bits_len(slave4.ARLEN),
        .slave4_ar_bits_size(slave4.ARSIZE),
        .slave4_ar_bits_burst(slave4.ARBURST),
        .slave4_ar_bits_lock(slave4.ARLOCK),
        .slave4_ar_bits_cache(slave4.ARCACHE),
        .slave4_ar_bits_prot(slave4.ARPROT),
        .slave4_ar_valid(slave4.ARVALID),
        .slave4_ar_ready(slave4.ARREADY),
        .slave4_r_bits_id(slave4.RID),
        .slave4_r_bits_data(slave4.RDATA),
        .slave4_r_bits_resp(slave4.RRESP),
        .slave4_r_bits_last(slave4.RLAST),
        .slave4_r_valid(slave4.RVALID),
        .slave4_r_ready(slave4.RREADY),
        .slave4_ar_bits_qos(slave4.ARQOS),
        .slave4_aw_bits_qos(slave4.AWQOS)        
      );


endmodule
/* verilator lint_on WIDTH */        

        
/* verilator lint_off WIDTH */        
module tb_AXI4XBar 
   (
   
   );

   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION master1;
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION master2;
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION slave1;
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION slave2;
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION slave3;
   AXI4_128_48_8_8_8_8_8_0_withQOS_noREGION slave4;
   logic  clock;
   logic  reset;


    AXI4XBar2x4 dut
      (
        .clock(clock),
        .reset(reset),
        .master1(master1),
        .master2(master2),
        .slave1(slave1),
        .slave2(slave2),
        .slave3(slave3),
        .slave4(slave4)        
      );


endmodule
/* verilator lint_on WIDTH */        
