
    // verilator lint_off DECLFILENAME
    // verilator lint_off UNUSED
    

interface AXI_4_53_1024_8_withQOS_noREGION;

   logic  ACLK;
   logic  ACLKEN;
   logic  ARESETn;
   logic [7:0] AWID;
   logic [52:0] AWADDR;
   logic [3:0] AWLEN;
   logic [2:0] AWSIZE;
   logic [1:0] AWBURST;
   logic [1:0] AWLOCK;
   logic [3:0] AWCACHE;
   logic [2:0] AWPROT;
   logic  AWVALID;
   logic  AWREADY;
   logic [7:0] WID;
   logic [1023:0] WDATA;
   logic [127:0] WSTRB;
   logic  WLAST;
   logic  WVALID;
   logic  WREADY;
   logic [7:0] BID;
   logic [1:0] BRESP;
   logic  BVALID;
   logic  BREADY;
   logic [7:0] ARID;
   logic [52:0] ARADDR;
   logic [3:0] ARLEN;
   logic [2:0] ARSIZE;
   logic [1:0] ARBURST;
   logic [1:0] ARLOCK;
   logic [3:0] ARCACHE;
   logic [2:0] ARPROT;
   logic  ARVALID;
   logic  ARREADY;
   logic [7:0] RID;
   logic [1023:0] RDATA;
   logic [1:0] RRESP;
   logic  RLAST;
   logic  RVALID;
   logic  RREADY;
   logic [7:0] AWUSER;
   logic [7:0] WUSER;
   logic [7:0] BUSER;
   logic [7:0] ARUSER;
   logic [7:0] RUSER;
   logic [3:0] ARQOS;
   logic [3:0] AWQOS;


    modport outward (
      input ACLK,
      input ACLKEN,
      input ARESETn,
      output AWID,
      output AWADDR,
      output AWLEN,
      output AWSIZE,
      output AWBURST,
      output AWLOCK,
      output AWCACHE,
      output AWPROT,
      output AWVALID,
      input AWREADY,
      output WID,
      output WDATA,
      output WSTRB,
      output WLAST,
      output WVALID,
      input WREADY,
      input BID,
      input BRESP,
      input BVALID,
      output BREADY,
      output ARID,
      output ARADDR,
      output ARLEN,
      output ARSIZE,
      output ARBURST,
      output ARLOCK,
      output ARCACHE,
      output ARPROT,
      output ARVALID,
      input ARREADY,
      input RID,
      input RDATA,
      input RRESP,
      input RLAST,
      input RVALID,
      output RREADY,
      output AWUSER,
      output WUSER,
      input BUSER,
      output ARUSER,
      input RUSER,
      output ARQOS,
      output AWQOS
    );           

    modport inward (
      output ACLK,
      output ACLKEN,
      output ARESETn,
      input AWID,
      input AWADDR,
      input AWLEN,
      input AWSIZE,
      input AWBURST,
      input AWLOCK,
      input AWCACHE,
      input AWPROT,
      input AWVALID,
      output AWREADY,
      input WID,
      input WDATA,
      input WSTRB,
      input WLAST,
      input WVALID,
      output WREADY,
      output BID,
      output BRESP,
      output BVALID,
      input BREADY,
      input ARID,
      input ARADDR,
      input ARLEN,
      input ARSIZE,
      input ARBURST,
      input ARLOCK,
      input ARCACHE,
      input ARPROT,
      input ARVALID,
      output ARREADY,
      output RID,
      output RDATA,
      output RRESP,
      output RLAST,
      output RVALID,
      input RREADY,
      input AWUSER,
      input WUSER,
      output BUSER,
      input ARUSER,
      output RUSER,
      input ARQOS,
      input AWQOS
    );           


endinterface
        
        
`timescale 1ps/1ps
module Specification_Architecture_Structure (
	Init0_Ar_Addr
,	Init0_Ar_Burst
,	Init0_Ar_Cache
,	Init0_Ar_Id
,	Init0_Ar_Len
,	Init0_Ar_Lock
,	Init0_Ar_Prot
,	Init0_Ar_Qos
,	Init0_Ar_Ready
,	Init0_Ar_Size
,	Init0_Ar_User
,	Init0_Ar_Valid
,	Init0_Aw_Addr
,	Init0_Aw_Burst
,	Init0_Aw_Cache
,	Init0_Aw_Id
,	Init0_Aw_Len
,	Init0_Aw_Lock
,	Init0_Aw_Prot
,	Init0_Aw_Qos
,	Init0_Aw_Ready
,	Init0_Aw_Size
,	Init0_Aw_User
,	Init0_Aw_Valid
,	Init0_B_Id
,	Init0_B_Ready
,	Init0_B_Resp
,	Init0_B_User
,	Init0_B_Valid
,	Init0_R_Data
,	Init0_R_Id
,	Init0_R_Last
,	Init0_R_Ready
,	Init0_R_Resp
,	Init0_R_User
,	Init0_R_Valid
,	Init0_W_Data
,	Init0_W_Id
,	Init0_W_Last
,	Init0_W_Ready
,	Init0_W_Strb
,	Init0_W_Valid
,	Init1_Ar_Addr
,	Init1_Ar_Burst
,	Init1_Ar_Cache
,	Init1_Ar_Id
,	Init1_Ar_Len
,	Init1_Ar_Lock
,	Init1_Ar_Prot
,	Init1_Ar_Qos
,	Init1_Ar_Ready
,	Init1_Ar_Size
,	Init1_Ar_User
,	Init1_Ar_Valid
,	Init1_Aw_Addr
,	Init1_Aw_Burst
,	Init1_Aw_Cache
,	Init1_Aw_Id
,	Init1_Aw_Len
,	Init1_Aw_Lock
,	Init1_Aw_Prot
,	Init1_Aw_Qos
,	Init1_Aw_Ready
,	Init1_Aw_Size
,	Init1_Aw_User
,	Init1_Aw_Valid
,	Init1_B_Id
,	Init1_B_Ready
,	Init1_B_Resp
,	Init1_B_User
,	Init1_B_Valid
,	Init1_R_Data
,	Init1_R_Id
,	Init1_R_Last
,	Init1_R_Ready
,	Init1_R_Resp
,	Init1_R_User
,	Init1_R_Valid
,	Init1_W_Data
,	Init1_W_Id
,	Init1_W_Last
,	Init1_W_Ready
,	Init1_W_Strb
,	Init1_W_Valid
,	Init10_Ar_Addr
,	Init10_Ar_Burst
,	Init10_Ar_Cache
,	Init10_Ar_Id
,	Init10_Ar_Len
,	Init10_Ar_Lock
,	Init10_Ar_Prot
,	Init10_Ar_Qos
,	Init10_Ar_Ready
,	Init10_Ar_Size
,	Init10_Ar_User
,	Init10_Ar_Valid
,	Init10_Aw_Addr
,	Init10_Aw_Burst
,	Init10_Aw_Cache
,	Init10_Aw_Id
,	Init10_Aw_Len
,	Init10_Aw_Lock
,	Init10_Aw_Prot
,	Init10_Aw_Qos
,	Init10_Aw_Ready
,	Init10_Aw_Size
,	Init10_Aw_User
,	Init10_Aw_Valid
,	Init10_B_Id
,	Init10_B_Ready
,	Init10_B_Resp
,	Init10_B_User
,	Init10_B_Valid
,	Init10_R_Data
,	Init10_R_Id
,	Init10_R_Last
,	Init10_R_Ready
,	Init10_R_Resp
,	Init10_R_User
,	Init10_R_Valid
,	Init10_W_Data
,	Init10_W_Id
,	Init10_W_Last
,	Init10_W_Ready
,	Init10_W_Strb
,	Init10_W_Valid
,	Init11_Ar_Addr
,	Init11_Ar_Burst
,	Init11_Ar_Cache
,	Init11_Ar_Id
,	Init11_Ar_Len
,	Init11_Ar_Lock
,	Init11_Ar_Prot
,	Init11_Ar_Qos
,	Init11_Ar_Ready
,	Init11_Ar_Size
,	Init11_Ar_User
,	Init11_Ar_Valid
,	Init11_Aw_Addr
,	Init11_Aw_Burst
,	Init11_Aw_Cache
,	Init11_Aw_Id
,	Init11_Aw_Len
,	Init11_Aw_Lock
,	Init11_Aw_Prot
,	Init11_Aw_Qos
,	Init11_Aw_Ready
,	Init11_Aw_Size
,	Init11_Aw_User
,	Init11_Aw_Valid
,	Init11_B_Id
,	Init11_B_Ready
,	Init11_B_Resp
,	Init11_B_User
,	Init11_B_Valid
,	Init11_R_Data
,	Init11_R_Id
,	Init11_R_Last
,	Init11_R_Ready
,	Init11_R_Resp
,	Init11_R_User
,	Init11_R_Valid
,	Init11_W_Data
,	Init11_W_Id
,	Init11_W_Last
,	Init11_W_Ready
,	Init11_W_Strb
,	Init11_W_Valid
,	Init2_Ar_Addr
,	Init2_Ar_Burst
,	Init2_Ar_Cache
,	Init2_Ar_Id
,	Init2_Ar_Len
,	Init2_Ar_Lock
,	Init2_Ar_Prot
,	Init2_Ar_Qos
,	Init2_Ar_Ready
,	Init2_Ar_Size
,	Init2_Ar_User
,	Init2_Ar_Valid
,	Init2_Aw_Addr
,	Init2_Aw_Burst
,	Init2_Aw_Cache
,	Init2_Aw_Id
,	Init2_Aw_Len
,	Init2_Aw_Lock
,	Init2_Aw_Prot
,	Init2_Aw_Qos
,	Init2_Aw_Ready
,	Init2_Aw_Size
,	Init2_Aw_User
,	Init2_Aw_Valid
,	Init2_B_Id
,	Init2_B_Ready
,	Init2_B_Resp
,	Init2_B_User
,	Init2_B_Valid
,	Init2_R_Data
,	Init2_R_Id
,	Init2_R_Last
,	Init2_R_Ready
,	Init2_R_Resp
,	Init2_R_User
,	Init2_R_Valid
,	Init2_W_Data
,	Init2_W_Id
,	Init2_W_Last
,	Init2_W_Ready
,	Init2_W_Strb
,	Init2_W_Valid
,	Init3_Ar_Addr
,	Init3_Ar_Burst
,	Init3_Ar_Cache
,	Init3_Ar_Id
,	Init3_Ar_Len
,	Init3_Ar_Lock
,	Init3_Ar_Prot
,	Init3_Ar_Qos
,	Init3_Ar_Ready
,	Init3_Ar_Size
,	Init3_Ar_User
,	Init3_Ar_Valid
,	Init3_Aw_Addr
,	Init3_Aw_Burst
,	Init3_Aw_Cache
,	Init3_Aw_Id
,	Init3_Aw_Len
,	Init3_Aw_Lock
,	Init3_Aw_Prot
,	Init3_Aw_Qos
,	Init3_Aw_Ready
,	Init3_Aw_Size
,	Init3_Aw_User
,	Init3_Aw_Valid
,	Init3_B_Id
,	Init3_B_Ready
,	Init3_B_Resp
,	Init3_B_User
,	Init3_B_Valid
,	Init3_R_Data
,	Init3_R_Id
,	Init3_R_Last
,	Init3_R_Ready
,	Init3_R_Resp
,	Init3_R_User
,	Init3_R_Valid
,	Init3_W_Data
,	Init3_W_Id
,	Init3_W_Last
,	Init3_W_Ready
,	Init3_W_Strb
,	Init3_W_Valid
,	Init4_Ar_Addr
,	Init4_Ar_Burst
,	Init4_Ar_Cache
,	Init4_Ar_Id
,	Init4_Ar_Len
,	Init4_Ar_Lock
,	Init4_Ar_Prot
,	Init4_Ar_Qos
,	Init4_Ar_Ready
,	Init4_Ar_Size
,	Init4_Ar_User
,	Init4_Ar_Valid
,	Init4_Aw_Addr
,	Init4_Aw_Burst
,	Init4_Aw_Cache
,	Init4_Aw_Id
,	Init4_Aw_Len
,	Init4_Aw_Lock
,	Init4_Aw_Prot
,	Init4_Aw_Qos
,	Init4_Aw_Ready
,	Init4_Aw_Size
,	Init4_Aw_User
,	Init4_Aw_Valid
,	Init4_B_Id
,	Init4_B_Ready
,	Init4_B_Resp
,	Init4_B_User
,	Init4_B_Valid
,	Init4_R_Data
,	Init4_R_Id
,	Init4_R_Last
,	Init4_R_Ready
,	Init4_R_Resp
,	Init4_R_User
,	Init4_R_Valid
,	Init4_W_Data
,	Init4_W_Id
,	Init4_W_Last
,	Init4_W_Ready
,	Init4_W_Strb
,	Init4_W_Valid
,	Init5_Ar_Addr
,	Init5_Ar_Burst
,	Init5_Ar_Cache
,	Init5_Ar_Id
,	Init5_Ar_Len
,	Init5_Ar_Lock
,	Init5_Ar_Prot
,	Init5_Ar_Qos
,	Init5_Ar_Ready
,	Init5_Ar_Size
,	Init5_Ar_User
,	Init5_Ar_Valid
,	Init5_Aw_Addr
,	Init5_Aw_Burst
,	Init5_Aw_Cache
,	Init5_Aw_Id
,	Init5_Aw_Len
,	Init5_Aw_Lock
,	Init5_Aw_Prot
,	Init5_Aw_Qos
,	Init5_Aw_Ready
,	Init5_Aw_Size
,	Init5_Aw_User
,	Init5_Aw_Valid
,	Init5_B_Id
,	Init5_B_Ready
,	Init5_B_Resp
,	Init5_B_User
,	Init5_B_Valid
,	Init5_R_Data
,	Init5_R_Id
,	Init5_R_Last
,	Init5_R_Ready
,	Init5_R_Resp
,	Init5_R_User
,	Init5_R_Valid
,	Init5_W_Data
,	Init5_W_Id
,	Init5_W_Last
,	Init5_W_Ready
,	Init5_W_Strb
,	Init5_W_Valid
,	Init6_Ar_Addr
,	Init6_Ar_Burst
,	Init6_Ar_Cache
,	Init6_Ar_Id
,	Init6_Ar_Len
,	Init6_Ar_Lock
,	Init6_Ar_Prot
,	Init6_Ar_Qos
,	Init6_Ar_Ready
,	Init6_Ar_Size
,	Init6_Ar_User
,	Init6_Ar_Valid
,	Init6_Aw_Addr
,	Init6_Aw_Burst
,	Init6_Aw_Cache
,	Init6_Aw_Id
,	Init6_Aw_Len
,	Init6_Aw_Lock
,	Init6_Aw_Prot
,	Init6_Aw_Qos
,	Init6_Aw_Ready
,	Init6_Aw_Size
,	Init6_Aw_User
,	Init6_Aw_Valid
,	Init6_B_Id
,	Init6_B_Ready
,	Init6_B_Resp
,	Init6_B_User
,	Init6_B_Valid
,	Init6_R_Data
,	Init6_R_Id
,	Init6_R_Last
,	Init6_R_Ready
,	Init6_R_Resp
,	Init6_R_User
,	Init6_R_Valid
,	Init6_W_Data
,	Init6_W_Id
,	Init6_W_Last
,	Init6_W_Ready
,	Init6_W_Strb
,	Init6_W_Valid
,	Init7_Ar_Addr
,	Init7_Ar_Burst
,	Init7_Ar_Cache
,	Init7_Ar_Id
,	Init7_Ar_Len
,	Init7_Ar_Lock
,	Init7_Ar_Prot
,	Init7_Ar_Qos
,	Init7_Ar_Ready
,	Init7_Ar_Size
,	Init7_Ar_User
,	Init7_Ar_Valid
,	Init7_Aw_Addr
,	Init7_Aw_Burst
,	Init7_Aw_Cache
,	Init7_Aw_Id
,	Init7_Aw_Len
,	Init7_Aw_Lock
,	Init7_Aw_Prot
,	Init7_Aw_Qos
,	Init7_Aw_Ready
,	Init7_Aw_Size
,	Init7_Aw_User
,	Init7_Aw_Valid
,	Init7_B_Id
,	Init7_B_Ready
,	Init7_B_Resp
,	Init7_B_User
,	Init7_B_Valid
,	Init7_R_Data
,	Init7_R_Id
,	Init7_R_Last
,	Init7_R_Ready
,	Init7_R_Resp
,	Init7_R_User
,	Init7_R_Valid
,	Init7_W_Data
,	Init7_W_Id
,	Init7_W_Last
,	Init7_W_Ready
,	Init7_W_Strb
,	Init7_W_Valid
,	Init8_Ar_Addr
,	Init8_Ar_Burst
,	Init8_Ar_Cache
,	Init8_Ar_Id
,	Init8_Ar_Len
,	Init8_Ar_Lock
,	Init8_Ar_Prot
,	Init8_Ar_Qos
,	Init8_Ar_Ready
,	Init8_Ar_Size
,	Init8_Ar_User
,	Init8_Ar_Valid
,	Init8_Aw_Addr
,	Init8_Aw_Burst
,	Init8_Aw_Cache
,	Init8_Aw_Id
,	Init8_Aw_Len
,	Init8_Aw_Lock
,	Init8_Aw_Prot
,	Init8_Aw_Qos
,	Init8_Aw_Ready
,	Init8_Aw_Size
,	Init8_Aw_User
,	Init8_Aw_Valid
,	Init8_B_Id
,	Init8_B_Ready
,	Init8_B_Resp
,	Init8_B_User
,	Init8_B_Valid
,	Init8_R_Data
,	Init8_R_Id
,	Init8_R_Last
,	Init8_R_Ready
,	Init8_R_Resp
,	Init8_R_User
,	Init8_R_Valid
,	Init8_W_Data
,	Init8_W_Id
,	Init8_W_Last
,	Init8_W_Ready
,	Init8_W_Strb
,	Init8_W_Valid
,	Init9_Ar_Addr
,	Init9_Ar_Burst
,	Init9_Ar_Cache
,	Init9_Ar_Id
,	Init9_Ar_Len
,	Init9_Ar_Lock
,	Init9_Ar_Prot
,	Init9_Ar_Qos
,	Init9_Ar_Ready
,	Init9_Ar_Size
,	Init9_Ar_User
,	Init9_Ar_Valid
,	Init9_Aw_Addr
,	Init9_Aw_Burst
,	Init9_Aw_Cache
,	Init9_Aw_Id
,	Init9_Aw_Len
,	Init9_Aw_Lock
,	Init9_Aw_Prot
,	Init9_Aw_Qos
,	Init9_Aw_Ready
,	Init9_Aw_Size
,	Init9_Aw_User
,	Init9_Aw_Valid
,	Init9_B_Id
,	Init9_B_Ready
,	Init9_B_Resp
,	Init9_B_User
,	Init9_B_Valid
,	Init9_R_Data
,	Init9_R_Id
,	Init9_R_Last
,	Init9_R_Ready
,	Init9_R_Resp
,	Init9_R_User
,	Init9_R_Valid
,	Init9_W_Data
,	Init9_W_Id
,	Init9_W_Last
,	Init9_W_Ready
,	Init9_W_Strb
,	Init9_W_Valid
,	Targ0_Ar_Addr
,	Targ0_Ar_Burst
,	Targ0_Ar_Cache
,	Targ0_Ar_Id
,	Targ0_Ar_Len
,	Targ0_Ar_Lock
,	Targ0_Ar_Prot
,	Targ0_Ar_Qos
,	Targ0_Ar_Ready
,	Targ0_Ar_Size
,	Targ0_Ar_User
,	Targ0_Ar_Valid
,	Targ0_Aw_Addr
,	Targ0_Aw_Burst
,	Targ0_Aw_Cache
,	Targ0_Aw_Id
,	Targ0_Aw_Len
,	Targ0_Aw_Lock
,	Targ0_Aw_Prot
,	Targ0_Aw_Qos
,	Targ0_Aw_Ready
,	Targ0_Aw_Size
,	Targ0_Aw_User
,	Targ0_Aw_Valid
,	Targ0_B_Id
,	Targ0_B_Ready
,	Targ0_B_Resp
,	Targ0_B_User
,	Targ0_B_Valid
,	Targ0_R_Data
,	Targ0_R_Id
,	Targ0_R_Last
,	Targ0_R_Ready
,	Targ0_R_Resp
,	Targ0_R_User
,	Targ0_R_Valid
,	Targ0_W_Data
,	Targ0_W_Id
,	Targ0_W_Last
,	Targ0_W_Ready
,	Targ0_W_Strb
,	Targ0_W_Valid
,	Targ1_Ar_Addr
,	Targ1_Ar_Burst
,	Targ1_Ar_Cache
,	Targ1_Ar_Id
,	Targ1_Ar_Len
,	Targ1_Ar_Lock
,	Targ1_Ar_Prot
,	Targ1_Ar_Qos
,	Targ1_Ar_Ready
,	Targ1_Ar_Size
,	Targ1_Ar_User
,	Targ1_Ar_Valid
,	Targ1_Aw_Addr
,	Targ1_Aw_Burst
,	Targ1_Aw_Cache
,	Targ1_Aw_Id
,	Targ1_Aw_Len
,	Targ1_Aw_Lock
,	Targ1_Aw_Prot
,	Targ1_Aw_Qos
,	Targ1_Aw_Ready
,	Targ1_Aw_Size
,	Targ1_Aw_User
,	Targ1_Aw_Valid
,	Targ1_B_Id
,	Targ1_B_Ready
,	Targ1_B_Resp
,	Targ1_B_User
,	Targ1_B_Valid
,	Targ1_R_Data
,	Targ1_R_Id
,	Targ1_R_Last
,	Targ1_R_Ready
,	Targ1_R_Resp
,	Targ1_R_User
,	Targ1_R_Valid
,	Targ1_W_Data
,	Targ1_W_Id
,	Targ1_W_Last
,	Targ1_W_Ready
,	Targ1_W_Strb
,	Targ1_W_Valid
,	Targ10_Ar_Addr
,	Targ10_Ar_Burst
,	Targ10_Ar_Cache
,	Targ10_Ar_Id
,	Targ10_Ar_Len
,	Targ10_Ar_Lock
,	Targ10_Ar_Prot
,	Targ10_Ar_Qos
,	Targ10_Ar_Ready
,	Targ10_Ar_Size
,	Targ10_Ar_User
,	Targ10_Ar_Valid
,	Targ10_Aw_Addr
,	Targ10_Aw_Burst
,	Targ10_Aw_Cache
,	Targ10_Aw_Id
,	Targ10_Aw_Len
,	Targ10_Aw_Lock
,	Targ10_Aw_Prot
,	Targ10_Aw_Qos
,	Targ10_Aw_Ready
,	Targ10_Aw_Size
,	Targ10_Aw_User
,	Targ10_Aw_Valid
,	Targ10_B_Id
,	Targ10_B_Ready
,	Targ10_B_Resp
,	Targ10_B_User
,	Targ10_B_Valid
,	Targ10_R_Data
,	Targ10_R_Id
,	Targ10_R_Last
,	Targ10_R_Ready
,	Targ10_R_Resp
,	Targ10_R_User
,	Targ10_R_Valid
,	Targ10_W_Data
,	Targ10_W_Id
,	Targ10_W_Last
,	Targ10_W_Ready
,	Targ10_W_Strb
,	Targ10_W_Valid
,	Targ11_Ar_Addr
,	Targ11_Ar_Burst
,	Targ11_Ar_Cache
,	Targ11_Ar_Id
,	Targ11_Ar_Len
,	Targ11_Ar_Lock
,	Targ11_Ar_Prot
,	Targ11_Ar_Qos
,	Targ11_Ar_Ready
,	Targ11_Ar_Size
,	Targ11_Ar_User
,	Targ11_Ar_Valid
,	Targ11_Aw_Addr
,	Targ11_Aw_Burst
,	Targ11_Aw_Cache
,	Targ11_Aw_Id
,	Targ11_Aw_Len
,	Targ11_Aw_Lock
,	Targ11_Aw_Prot
,	Targ11_Aw_Qos
,	Targ11_Aw_Ready
,	Targ11_Aw_Size
,	Targ11_Aw_User
,	Targ11_Aw_Valid
,	Targ11_B_Id
,	Targ11_B_Ready
,	Targ11_B_Resp
,	Targ11_B_User
,	Targ11_B_Valid
,	Targ11_R_Data
,	Targ11_R_Id
,	Targ11_R_Last
,	Targ11_R_Ready
,	Targ11_R_Resp
,	Targ11_R_User
,	Targ11_R_Valid
,	Targ11_W_Data
,	Targ11_W_Id
,	Targ11_W_Last
,	Targ11_W_Ready
,	Targ11_W_Strb
,	Targ11_W_Valid
,	Targ2_Ar_Addr
,	Targ2_Ar_Burst
,	Targ2_Ar_Cache
,	Targ2_Ar_Id
,	Targ2_Ar_Len
,	Targ2_Ar_Lock
,	Targ2_Ar_Prot
,	Targ2_Ar_Qos
,	Targ2_Ar_Ready
,	Targ2_Ar_Size
,	Targ2_Ar_User
,	Targ2_Ar_Valid
,	Targ2_Aw_Addr
,	Targ2_Aw_Burst
,	Targ2_Aw_Cache
,	Targ2_Aw_Id
,	Targ2_Aw_Len
,	Targ2_Aw_Lock
,	Targ2_Aw_Prot
,	Targ2_Aw_Qos
,	Targ2_Aw_Ready
,	Targ2_Aw_Size
,	Targ2_Aw_User
,	Targ2_Aw_Valid
,	Targ2_B_Id
,	Targ2_B_Ready
,	Targ2_B_Resp
,	Targ2_B_User
,	Targ2_B_Valid
,	Targ2_R_Data
,	Targ2_R_Id
,	Targ2_R_Last
,	Targ2_R_Ready
,	Targ2_R_Resp
,	Targ2_R_User
,	Targ2_R_Valid
,	Targ2_W_Data
,	Targ2_W_Id
,	Targ2_W_Last
,	Targ2_W_Ready
,	Targ2_W_Strb
,	Targ2_W_Valid
,	Targ3_Ar_Addr
,	Targ3_Ar_Burst
,	Targ3_Ar_Cache
,	Targ3_Ar_Id
,	Targ3_Ar_Len
,	Targ3_Ar_Lock
,	Targ3_Ar_Prot
,	Targ3_Ar_Qos
,	Targ3_Ar_Ready
,	Targ3_Ar_Size
,	Targ3_Ar_User
,	Targ3_Ar_Valid
,	Targ3_Aw_Addr
,	Targ3_Aw_Burst
,	Targ3_Aw_Cache
,	Targ3_Aw_Id
,	Targ3_Aw_Len
,	Targ3_Aw_Lock
,	Targ3_Aw_Prot
,	Targ3_Aw_Qos
,	Targ3_Aw_Ready
,	Targ3_Aw_Size
,	Targ3_Aw_User
,	Targ3_Aw_Valid
,	Targ3_B_Id
,	Targ3_B_Ready
,	Targ3_B_Resp
,	Targ3_B_User
,	Targ3_B_Valid
,	Targ3_R_Data
,	Targ3_R_Id
,	Targ3_R_Last
,	Targ3_R_Ready
,	Targ3_R_Resp
,	Targ3_R_User
,	Targ3_R_Valid
,	Targ3_W_Data
,	Targ3_W_Id
,	Targ3_W_Last
,	Targ3_W_Ready
,	Targ3_W_Strb
,	Targ3_W_Valid
,	Targ4_Ar_Addr
,	Targ4_Ar_Burst
,	Targ4_Ar_Cache
,	Targ4_Ar_Id
,	Targ4_Ar_Len
,	Targ4_Ar_Lock
,	Targ4_Ar_Prot
,	Targ4_Ar_Qos
,	Targ4_Ar_Ready
,	Targ4_Ar_Size
,	Targ4_Ar_User
,	Targ4_Ar_Valid
,	Targ4_Aw_Addr
,	Targ4_Aw_Burst
,	Targ4_Aw_Cache
,	Targ4_Aw_Id
,	Targ4_Aw_Len
,	Targ4_Aw_Lock
,	Targ4_Aw_Prot
,	Targ4_Aw_Qos
,	Targ4_Aw_Ready
,	Targ4_Aw_Size
,	Targ4_Aw_User
,	Targ4_Aw_Valid
,	Targ4_B_Id
,	Targ4_B_Ready
,	Targ4_B_Resp
,	Targ4_B_User
,	Targ4_B_Valid
,	Targ4_R_Data
,	Targ4_R_Id
,	Targ4_R_Last
,	Targ4_R_Ready
,	Targ4_R_Resp
,	Targ4_R_User
,	Targ4_R_Valid
,	Targ4_W_Data
,	Targ4_W_Id
,	Targ4_W_Last
,	Targ4_W_Ready
,	Targ4_W_Strb
,	Targ4_W_Valid
,	Targ5_Ar_Addr
,	Targ5_Ar_Burst
,	Targ5_Ar_Cache
,	Targ5_Ar_Id
,	Targ5_Ar_Len
,	Targ5_Ar_Lock
,	Targ5_Ar_Prot
,	Targ5_Ar_Qos
,	Targ5_Ar_Ready
,	Targ5_Ar_Size
,	Targ5_Ar_User
,	Targ5_Ar_Valid
,	Targ5_Aw_Addr
,	Targ5_Aw_Burst
,	Targ5_Aw_Cache
,	Targ5_Aw_Id
,	Targ5_Aw_Len
,	Targ5_Aw_Lock
,	Targ5_Aw_Prot
,	Targ5_Aw_Qos
,	Targ5_Aw_Ready
,	Targ5_Aw_Size
,	Targ5_Aw_User
,	Targ5_Aw_Valid
,	Targ5_B_Id
,	Targ5_B_Ready
,	Targ5_B_Resp
,	Targ5_B_User
,	Targ5_B_Valid
,	Targ5_R_Data
,	Targ5_R_Id
,	Targ5_R_Last
,	Targ5_R_Ready
,	Targ5_R_Resp
,	Targ5_R_User
,	Targ5_R_Valid
,	Targ5_W_Data
,	Targ5_W_Id
,	Targ5_W_Last
,	Targ5_W_Ready
,	Targ5_W_Strb
,	Targ5_W_Valid
,	Targ6_Ar_Addr
,	Targ6_Ar_Burst
,	Targ6_Ar_Cache
,	Targ6_Ar_Id
,	Targ6_Ar_Len
,	Targ6_Ar_Lock
,	Targ6_Ar_Prot
,	Targ6_Ar_Qos
,	Targ6_Ar_Ready
,	Targ6_Ar_Size
,	Targ6_Ar_User
,	Targ6_Ar_Valid
,	Targ6_Aw_Addr
,	Targ6_Aw_Burst
,	Targ6_Aw_Cache
,	Targ6_Aw_Id
,	Targ6_Aw_Len
,	Targ6_Aw_Lock
,	Targ6_Aw_Prot
,	Targ6_Aw_Qos
,	Targ6_Aw_Ready
,	Targ6_Aw_Size
,	Targ6_Aw_User
,	Targ6_Aw_Valid
,	Targ6_B_Id
,	Targ6_B_Ready
,	Targ6_B_Resp
,	Targ6_B_User
,	Targ6_B_Valid
,	Targ6_R_Data
,	Targ6_R_Id
,	Targ6_R_Last
,	Targ6_R_Ready
,	Targ6_R_Resp
,	Targ6_R_User
,	Targ6_R_Valid
,	Targ6_W_Data
,	Targ6_W_Id
,	Targ6_W_Last
,	Targ6_W_Ready
,	Targ6_W_Strb
,	Targ6_W_Valid
,	Targ7_Ar_Addr
,	Targ7_Ar_Burst
,	Targ7_Ar_Cache
,	Targ7_Ar_Id
,	Targ7_Ar_Len
,	Targ7_Ar_Lock
,	Targ7_Ar_Prot
,	Targ7_Ar_Qos
,	Targ7_Ar_Ready
,	Targ7_Ar_Size
,	Targ7_Ar_User
,	Targ7_Ar_Valid
,	Targ7_Aw_Addr
,	Targ7_Aw_Burst
,	Targ7_Aw_Cache
,	Targ7_Aw_Id
,	Targ7_Aw_Len
,	Targ7_Aw_Lock
,	Targ7_Aw_Prot
,	Targ7_Aw_Qos
,	Targ7_Aw_Ready
,	Targ7_Aw_Size
,	Targ7_Aw_User
,	Targ7_Aw_Valid
,	Targ7_B_Id
,	Targ7_B_Ready
,	Targ7_B_Resp
,	Targ7_B_User
,	Targ7_B_Valid
,	Targ7_R_Data
,	Targ7_R_Id
,	Targ7_R_Last
,	Targ7_R_Ready
,	Targ7_R_Resp
,	Targ7_R_User
,	Targ7_R_Valid
,	Targ7_W_Data
,	Targ7_W_Id
,	Targ7_W_Last
,	Targ7_W_Ready
,	Targ7_W_Strb
,	Targ7_W_Valid
,	Targ8_Ar_Addr
,	Targ8_Ar_Burst
,	Targ8_Ar_Cache
,	Targ8_Ar_Id
,	Targ8_Ar_Len
,	Targ8_Ar_Lock
,	Targ8_Ar_Prot
,	Targ8_Ar_Qos
,	Targ8_Ar_Ready
,	Targ8_Ar_Size
,	Targ8_Ar_User
,	Targ8_Ar_Valid
,	Targ8_Aw_Addr
,	Targ8_Aw_Burst
,	Targ8_Aw_Cache
,	Targ8_Aw_Id
,	Targ8_Aw_Len
,	Targ8_Aw_Lock
,	Targ8_Aw_Prot
,	Targ8_Aw_Qos
,	Targ8_Aw_Ready
,	Targ8_Aw_Size
,	Targ8_Aw_User
,	Targ8_Aw_Valid
,	Targ8_B_Id
,	Targ8_B_Ready
,	Targ8_B_Resp
,	Targ8_B_User
,	Targ8_B_Valid
,	Targ8_R_Data
,	Targ8_R_Id
,	Targ8_R_Last
,	Targ8_R_Ready
,	Targ8_R_Resp
,	Targ8_R_User
,	Targ8_R_Valid
,	Targ8_W_Data
,	Targ8_W_Id
,	Targ8_W_Last
,	Targ8_W_Ready
,	Targ8_W_Strb
,	Targ8_W_Valid
,	Targ9_Ar_Addr
,	Targ9_Ar_Burst
,	Targ9_Ar_Cache
,	Targ9_Ar_Id
,	Targ9_Ar_Len
,	Targ9_Ar_Lock
,	Targ9_Ar_Prot
,	Targ9_Ar_Qos
,	Targ9_Ar_Ready
,	Targ9_Ar_Size
,	Targ9_Ar_User
,	Targ9_Ar_Valid
,	Targ9_Aw_Addr
,	Targ9_Aw_Burst
,	Targ9_Aw_Cache
,	Targ9_Aw_Id
,	Targ9_Aw_Len
,	Targ9_Aw_Lock
,	Targ9_Aw_Prot
,	Targ9_Aw_Qos
,	Targ9_Aw_Ready
,	Targ9_Aw_Size
,	Targ9_Aw_User
,	Targ9_Aw_Valid
,	Targ9_B_Id
,	Targ9_B_Ready
,	Targ9_B_Resp
,	Targ9_B_User
,	Targ9_B_Valid
,	Targ9_R_Data
,	Targ9_R_Id
,	Targ9_R_Last
,	Targ9_R_Ready
,	Targ9_R_Resp
,	Targ9_R_User
,	Targ9_R_Valid
,	Targ9_W_Data
,	Targ9_W_Id
,	Targ9_W_Last
,	Targ9_W_Ready
,	Targ9_W_Strb
,	Targ9_W_Valid
,	noc_arstn
,	node0_aclk
,	node10_aclk
,	node11_aclk
,	node1_aclk
,	node2_aclk
,	node3_aclk
,	node4_aclk
,	node5_aclk
,	node6_aclk
,	node7_aclk
,	node8_aclk
,	node9_aclk
,	tm
);
	input  [52:0]   Init0_Ar_Addr   ;
	input  [1:0]    Init0_Ar_Burst  ;
	input  [3:0]    Init0_Ar_Cache  ;
	input  [7:0]    Init0_Ar_Id     ;
	input  [7:0]    Init0_Ar_Len    ;
	input  [1:0]    Init0_Ar_Lock   ;
	input  [2:0]    Init0_Ar_Prot   ;
	input  [3:0]    Init0_Ar_Qos    ;
	output          Init0_Ar_Ready  ;
	input  [2:0]    Init0_Ar_Size   ;
	input  [7:0]    Init0_Ar_User   ;
	input           Init0_Ar_Valid  ;
	input  [52:0]   Init0_Aw_Addr   ;
	input  [1:0]    Init0_Aw_Burst  ;
	input  [3:0]    Init0_Aw_Cache  ;
	input  [7:0]    Init0_Aw_Id     ;
	input  [7:0]    Init0_Aw_Len    ;
	input  [1:0]    Init0_Aw_Lock   ;
	input  [2:0]    Init0_Aw_Prot   ;
	input  [3:0]    Init0_Aw_Qos    ;
	output          Init0_Aw_Ready  ;
	input  [2:0]    Init0_Aw_Size   ;
	input  [7:0]    Init0_Aw_User   ;
	input           Init0_Aw_Valid  ;
	output [7:0]    Init0_B_Id      ;
	input           Init0_B_Ready   ;
	output [1:0]    Init0_B_Resp    ;
	output [7:0]    Init0_B_User    ;
	output          Init0_B_Valid   ;
	output [1023:0] Init0_R_Data    ;
	output [7:0]    Init0_R_Id      ;
	output          Init0_R_Last    ;
	input           Init0_R_Ready   ;
	output [1:0]    Init0_R_Resp    ;
	output [7:0]    Init0_R_User    ;
	output          Init0_R_Valid   ;
	input  [1023:0] Init0_W_Data    ;
	input  [7:0]    Init0_W_Id      ;
	input           Init0_W_Last    ;
	output          Init0_W_Ready   ;
	input  [127:0]  Init0_W_Strb    ;
	input           Init0_W_Valid   ;
	input  [52:0]   Init1_Ar_Addr   ;
	input  [1:0]    Init1_Ar_Burst  ;
	input  [3:0]    Init1_Ar_Cache  ;
	input  [7:0]    Init1_Ar_Id     ;
	input  [7:0]    Init1_Ar_Len    ;
	input  [1:0]    Init1_Ar_Lock   ;
	input  [2:0]    Init1_Ar_Prot   ;
	input  [3:0]    Init1_Ar_Qos    ;
	output          Init1_Ar_Ready  ;
	input  [2:0]    Init1_Ar_Size   ;
	input  [7:0]    Init1_Ar_User   ;
	input           Init1_Ar_Valid  ;
	input  [52:0]   Init1_Aw_Addr   ;
	input  [1:0]    Init1_Aw_Burst  ;
	input  [3:0]    Init1_Aw_Cache  ;
	input  [7:0]    Init1_Aw_Id     ;
	input  [7:0]    Init1_Aw_Len    ;
	input  [1:0]    Init1_Aw_Lock   ;
	input  [2:0]    Init1_Aw_Prot   ;
	input  [3:0]    Init1_Aw_Qos    ;
	output          Init1_Aw_Ready  ;
	input  [2:0]    Init1_Aw_Size   ;
	input  [7:0]    Init1_Aw_User   ;
	input           Init1_Aw_Valid  ;
	output [7:0]    Init1_B_Id      ;
	input           Init1_B_Ready   ;
	output [1:0]    Init1_B_Resp    ;
	output [7:0]    Init1_B_User    ;
	output          Init1_B_Valid   ;
	output [1023:0] Init1_R_Data    ;
	output [7:0]    Init1_R_Id      ;
	output          Init1_R_Last    ;
	input           Init1_R_Ready   ;
	output [1:0]    Init1_R_Resp    ;
	output [7:0]    Init1_R_User    ;
	output          Init1_R_Valid   ;
	input  [1023:0] Init1_W_Data    ;
	input  [7:0]    Init1_W_Id      ;
	input           Init1_W_Last    ;
	output          Init1_W_Ready   ;
	input  [127:0]  Init1_W_Strb    ;
	input           Init1_W_Valid   ;
	input  [52:0]   Init10_Ar_Addr  ;
	input  [1:0]    Init10_Ar_Burst ;
	input  [3:0]    Init10_Ar_Cache ;
	input  [7:0]    Init10_Ar_Id    ;
	input  [7:0]    Init10_Ar_Len   ;
	input  [1:0]    Init10_Ar_Lock  ;
	input  [2:0]    Init10_Ar_Prot  ;
	input  [3:0]    Init10_Ar_Qos   ;
	output          Init10_Ar_Ready ;
	input  [2:0]    Init10_Ar_Size  ;
	input  [7:0]    Init10_Ar_User  ;
	input           Init10_Ar_Valid ;
	input  [52:0]   Init10_Aw_Addr  ;
	input  [1:0]    Init10_Aw_Burst ;
	input  [3:0]    Init10_Aw_Cache ;
	input  [7:0]    Init10_Aw_Id    ;
	input  [7:0]    Init10_Aw_Len   ;
	input  [1:0]    Init10_Aw_Lock  ;
	input  [2:0]    Init10_Aw_Prot  ;
	input  [3:0]    Init10_Aw_Qos   ;
	output          Init10_Aw_Ready ;
	input  [2:0]    Init10_Aw_Size  ;
	input  [7:0]    Init10_Aw_User  ;
	input           Init10_Aw_Valid ;
	output [7:0]    Init10_B_Id     ;
	input           Init10_B_Ready  ;
	output [1:0]    Init10_B_Resp   ;
	output [7:0]    Init10_B_User   ;
	output          Init10_B_Valid  ;
	output [1023:0] Init10_R_Data   ;
	output [7:0]    Init10_R_Id     ;
	output          Init10_R_Last   ;
	input           Init10_R_Ready  ;
	output [1:0]    Init10_R_Resp   ;
	output [7:0]    Init10_R_User   ;
	output          Init10_R_Valid  ;
	input  [1023:0] Init10_W_Data   ;
	input  [7:0]    Init10_W_Id     ;
	input           Init10_W_Last   ;
	output          Init10_W_Ready  ;
	input  [127:0]  Init10_W_Strb   ;
	input           Init10_W_Valid  ;
	input  [52:0]   Init11_Ar_Addr  ;
	input  [1:0]    Init11_Ar_Burst ;
	input  [3:0]    Init11_Ar_Cache ;
	input  [7:0]    Init11_Ar_Id    ;
	input  [7:0]    Init11_Ar_Len   ;
	input  [1:0]    Init11_Ar_Lock  ;
	input  [2:0]    Init11_Ar_Prot  ;
	input  [3:0]    Init11_Ar_Qos   ;
	output          Init11_Ar_Ready ;
	input  [2:0]    Init11_Ar_Size  ;
	input  [7:0]    Init11_Ar_User  ;
	input           Init11_Ar_Valid ;
	input  [52:0]   Init11_Aw_Addr  ;
	input  [1:0]    Init11_Aw_Burst ;
	input  [3:0]    Init11_Aw_Cache ;
	input  [7:0]    Init11_Aw_Id    ;
	input  [7:0]    Init11_Aw_Len   ;
	input  [1:0]    Init11_Aw_Lock  ;
	input  [2:0]    Init11_Aw_Prot  ;
	input  [3:0]    Init11_Aw_Qos   ;
	output          Init11_Aw_Ready ;
	input  [2:0]    Init11_Aw_Size  ;
	input  [7:0]    Init11_Aw_User  ;
	input           Init11_Aw_Valid ;
	output [7:0]    Init11_B_Id     ;
	input           Init11_B_Ready  ;
	output [1:0]    Init11_B_Resp   ;
	output [7:0]    Init11_B_User   ;
	output          Init11_B_Valid  ;
	output [1023:0] Init11_R_Data   ;
	output [7:0]    Init11_R_Id     ;
	output          Init11_R_Last   ;
	input           Init11_R_Ready  ;
	output [1:0]    Init11_R_Resp   ;
	output [7:0]    Init11_R_User   ;
	output          Init11_R_Valid  ;
	input  [1023:0] Init11_W_Data   ;
	input  [7:0]    Init11_W_Id     ;
	input           Init11_W_Last   ;
	output          Init11_W_Ready  ;
	input  [127:0]  Init11_W_Strb   ;
	input           Init11_W_Valid  ;
	input  [52:0]   Init2_Ar_Addr   ;
	input  [1:0]    Init2_Ar_Burst  ;
	input  [3:0]    Init2_Ar_Cache  ;
	input  [7:0]    Init2_Ar_Id     ;
	input  [7:0]    Init2_Ar_Len    ;
	input  [1:0]    Init2_Ar_Lock   ;
	input  [2:0]    Init2_Ar_Prot   ;
	input  [3:0]    Init2_Ar_Qos    ;
	output          Init2_Ar_Ready  ;
	input  [2:0]    Init2_Ar_Size   ;
	input  [7:0]    Init2_Ar_User   ;
	input           Init2_Ar_Valid  ;
	input  [52:0]   Init2_Aw_Addr   ;
	input  [1:0]    Init2_Aw_Burst  ;
	input  [3:0]    Init2_Aw_Cache  ;
	input  [7:0]    Init2_Aw_Id     ;
	input  [7:0]    Init2_Aw_Len    ;
	input  [1:0]    Init2_Aw_Lock   ;
	input  [2:0]    Init2_Aw_Prot   ;
	input  [3:0]    Init2_Aw_Qos    ;
	output          Init2_Aw_Ready  ;
	input  [2:0]    Init2_Aw_Size   ;
	input  [7:0]    Init2_Aw_User   ;
	input           Init2_Aw_Valid  ;
	output [7:0]    Init2_B_Id      ;
	input           Init2_B_Ready   ;
	output [1:0]    Init2_B_Resp    ;
	output [7:0]    Init2_B_User    ;
	output          Init2_B_Valid   ;
	output [1023:0] Init2_R_Data    ;
	output [7:0]    Init2_R_Id      ;
	output          Init2_R_Last    ;
	input           Init2_R_Ready   ;
	output [1:0]    Init2_R_Resp    ;
	output [7:0]    Init2_R_User    ;
	output          Init2_R_Valid   ;
	input  [1023:0] Init2_W_Data    ;
	input  [7:0]    Init2_W_Id      ;
	input           Init2_W_Last    ;
	output          Init2_W_Ready   ;
	input  [127:0]  Init2_W_Strb    ;
	input           Init2_W_Valid   ;
	input  [52:0]   Init3_Ar_Addr   ;
	input  [1:0]    Init3_Ar_Burst  ;
	input  [3:0]    Init3_Ar_Cache  ;
	input  [7:0]    Init3_Ar_Id     ;
	input  [7:0]    Init3_Ar_Len    ;
	input  [1:0]    Init3_Ar_Lock   ;
	input  [2:0]    Init3_Ar_Prot   ;
	input  [3:0]    Init3_Ar_Qos    ;
	output          Init3_Ar_Ready  ;
	input  [2:0]    Init3_Ar_Size   ;
	input  [7:0]    Init3_Ar_User   ;
	input           Init3_Ar_Valid  ;
	input  [52:0]   Init3_Aw_Addr   ;
	input  [1:0]    Init3_Aw_Burst  ;
	input  [3:0]    Init3_Aw_Cache  ;
	input  [7:0]    Init3_Aw_Id     ;
	input  [7:0]    Init3_Aw_Len    ;
	input  [1:0]    Init3_Aw_Lock   ;
	input  [2:0]    Init3_Aw_Prot   ;
	input  [3:0]    Init3_Aw_Qos    ;
	output          Init3_Aw_Ready  ;
	input  [2:0]    Init3_Aw_Size   ;
	input  [7:0]    Init3_Aw_User   ;
	input           Init3_Aw_Valid  ;
	output [7:0]    Init3_B_Id      ;
	input           Init3_B_Ready   ;
	output [1:0]    Init3_B_Resp    ;
	output [7:0]    Init3_B_User    ;
	output          Init3_B_Valid   ;
	output [1023:0] Init3_R_Data    ;
	output [7:0]    Init3_R_Id      ;
	output          Init3_R_Last    ;
	input           Init3_R_Ready   ;
	output [1:0]    Init3_R_Resp    ;
	output [7:0]    Init3_R_User    ;
	output          Init3_R_Valid   ;
	input  [1023:0] Init3_W_Data    ;
	input  [7:0]    Init3_W_Id      ;
	input           Init3_W_Last    ;
	output          Init3_W_Ready   ;
	input  [127:0]  Init3_W_Strb    ;
	input           Init3_W_Valid   ;
	input  [52:0]   Init4_Ar_Addr   ;
	input  [1:0]    Init4_Ar_Burst  ;
	input  [3:0]    Init4_Ar_Cache  ;
	input  [7:0]    Init4_Ar_Id     ;
	input  [7:0]    Init4_Ar_Len    ;
	input  [1:0]    Init4_Ar_Lock   ;
	input  [2:0]    Init4_Ar_Prot   ;
	input  [3:0]    Init4_Ar_Qos    ;
	output          Init4_Ar_Ready  ;
	input  [2:0]    Init4_Ar_Size   ;
	input  [7:0]    Init4_Ar_User   ;
	input           Init4_Ar_Valid  ;
	input  [52:0]   Init4_Aw_Addr   ;
	input  [1:0]    Init4_Aw_Burst  ;
	input  [3:0]    Init4_Aw_Cache  ;
	input  [7:0]    Init4_Aw_Id     ;
	input  [7:0]    Init4_Aw_Len    ;
	input  [1:0]    Init4_Aw_Lock   ;
	input  [2:0]    Init4_Aw_Prot   ;
	input  [3:0]    Init4_Aw_Qos    ;
	output          Init4_Aw_Ready  ;
	input  [2:0]    Init4_Aw_Size   ;
	input  [7:0]    Init4_Aw_User   ;
	input           Init4_Aw_Valid  ;
	output [7:0]    Init4_B_Id      ;
	input           Init4_B_Ready   ;
	output [1:0]    Init4_B_Resp    ;
	output [7:0]    Init4_B_User    ;
	output          Init4_B_Valid   ;
	output [1023:0] Init4_R_Data    ;
	output [7:0]    Init4_R_Id      ;
	output          Init4_R_Last    ;
	input           Init4_R_Ready   ;
	output [1:0]    Init4_R_Resp    ;
	output [7:0]    Init4_R_User    ;
	output          Init4_R_Valid   ;
	input  [1023:0] Init4_W_Data    ;
	input  [7:0]    Init4_W_Id      ;
	input           Init4_W_Last    ;
	output          Init4_W_Ready   ;
	input  [127:0]  Init4_W_Strb    ;
	input           Init4_W_Valid   ;
	input  [52:0]   Init5_Ar_Addr   ;
	input  [1:0]    Init5_Ar_Burst  ;
	input  [3:0]    Init5_Ar_Cache  ;
	input  [7:0]    Init5_Ar_Id     ;
	input  [7:0]    Init5_Ar_Len    ;
	input  [1:0]    Init5_Ar_Lock   ;
	input  [2:0]    Init5_Ar_Prot   ;
	input  [3:0]    Init5_Ar_Qos    ;
	output          Init5_Ar_Ready  ;
	input  [2:0]    Init5_Ar_Size   ;
	input  [7:0]    Init5_Ar_User   ;
	input           Init5_Ar_Valid  ;
	input  [52:0]   Init5_Aw_Addr   ;
	input  [1:0]    Init5_Aw_Burst  ;
	input  [3:0]    Init5_Aw_Cache  ;
	input  [7:0]    Init5_Aw_Id     ;
	input  [7:0]    Init5_Aw_Len    ;
	input  [1:0]    Init5_Aw_Lock   ;
	input  [2:0]    Init5_Aw_Prot   ;
	input  [3:0]    Init5_Aw_Qos    ;
	output          Init5_Aw_Ready  ;
	input  [2:0]    Init5_Aw_Size   ;
	input  [7:0]    Init5_Aw_User   ;
	input           Init5_Aw_Valid  ;
	output [7:0]    Init5_B_Id      ;
	input           Init5_B_Ready   ;
	output [1:0]    Init5_B_Resp    ;
	output [7:0]    Init5_B_User    ;
	output          Init5_B_Valid   ;
	output [1023:0] Init5_R_Data    ;
	output [7:0]    Init5_R_Id      ;
	output          Init5_R_Last    ;
	input           Init5_R_Ready   ;
	output [1:0]    Init5_R_Resp    ;
	output [7:0]    Init5_R_User    ;
	output          Init5_R_Valid   ;
	input  [1023:0] Init5_W_Data    ;
	input  [7:0]    Init5_W_Id      ;
	input           Init5_W_Last    ;
	output          Init5_W_Ready   ;
	input  [127:0]  Init5_W_Strb    ;
	input           Init5_W_Valid   ;
	input  [52:0]   Init6_Ar_Addr   ;
	input  [1:0]    Init6_Ar_Burst  ;
	input  [3:0]    Init6_Ar_Cache  ;
	input  [7:0]    Init6_Ar_Id     ;
	input  [7:0]    Init6_Ar_Len    ;
	input  [1:0]    Init6_Ar_Lock   ;
	input  [2:0]    Init6_Ar_Prot   ;
	input  [3:0]    Init6_Ar_Qos    ;
	output          Init6_Ar_Ready  ;
	input  [2:0]    Init6_Ar_Size   ;
	input  [7:0]    Init6_Ar_User   ;
	input           Init6_Ar_Valid  ;
	input  [52:0]   Init6_Aw_Addr   ;
	input  [1:0]    Init6_Aw_Burst  ;
	input  [3:0]    Init6_Aw_Cache  ;
	input  [7:0]    Init6_Aw_Id     ;
	input  [7:0]    Init6_Aw_Len    ;
	input  [1:0]    Init6_Aw_Lock   ;
	input  [2:0]    Init6_Aw_Prot   ;
	input  [3:0]    Init6_Aw_Qos    ;
	output          Init6_Aw_Ready  ;
	input  [2:0]    Init6_Aw_Size   ;
	input  [7:0]    Init6_Aw_User   ;
	input           Init6_Aw_Valid  ;
	output [7:0]    Init6_B_Id      ;
	input           Init6_B_Ready   ;
	output [1:0]    Init6_B_Resp    ;
	output [7:0]    Init6_B_User    ;
	output          Init6_B_Valid   ;
	output [1023:0] Init6_R_Data    ;
	output [7:0]    Init6_R_Id      ;
	output          Init6_R_Last    ;
	input           Init6_R_Ready   ;
	output [1:0]    Init6_R_Resp    ;
	output [7:0]    Init6_R_User    ;
	output          Init6_R_Valid   ;
	input  [1023:0] Init6_W_Data    ;
	input  [7:0]    Init6_W_Id      ;
	input           Init6_W_Last    ;
	output          Init6_W_Ready   ;
	input  [127:0]  Init6_W_Strb    ;
	input           Init6_W_Valid   ;
	input  [52:0]   Init7_Ar_Addr   ;
	input  [1:0]    Init7_Ar_Burst  ;
	input  [3:0]    Init7_Ar_Cache  ;
	input  [7:0]    Init7_Ar_Id     ;
	input  [7:0]    Init7_Ar_Len    ;
	input  [1:0]    Init7_Ar_Lock   ;
	input  [2:0]    Init7_Ar_Prot   ;
	input  [3:0]    Init7_Ar_Qos    ;
	output          Init7_Ar_Ready  ;
	input  [2:0]    Init7_Ar_Size   ;
	input  [7:0]    Init7_Ar_User   ;
	input           Init7_Ar_Valid  ;
	input  [52:0]   Init7_Aw_Addr   ;
	input  [1:0]    Init7_Aw_Burst  ;
	input  [3:0]    Init7_Aw_Cache  ;
	input  [7:0]    Init7_Aw_Id     ;
	input  [7:0]    Init7_Aw_Len    ;
	input  [1:0]    Init7_Aw_Lock   ;
	input  [2:0]    Init7_Aw_Prot   ;
	input  [3:0]    Init7_Aw_Qos    ;
	output          Init7_Aw_Ready  ;
	input  [2:0]    Init7_Aw_Size   ;
	input  [7:0]    Init7_Aw_User   ;
	input           Init7_Aw_Valid  ;
	output [7:0]    Init7_B_Id      ;
	input           Init7_B_Ready   ;
	output [1:0]    Init7_B_Resp    ;
	output [7:0]    Init7_B_User    ;
	output          Init7_B_Valid   ;
	output [1023:0] Init7_R_Data    ;
	output [7:0]    Init7_R_Id      ;
	output          Init7_R_Last    ;
	input           Init7_R_Ready   ;
	output [1:0]    Init7_R_Resp    ;
	output [7:0]    Init7_R_User    ;
	output          Init7_R_Valid   ;
	input  [1023:0] Init7_W_Data    ;
	input  [7:0]    Init7_W_Id      ;
	input           Init7_W_Last    ;
	output          Init7_W_Ready   ;
	input  [127:0]  Init7_W_Strb    ;
	input           Init7_W_Valid   ;
	input  [52:0]   Init8_Ar_Addr   ;
	input  [1:0]    Init8_Ar_Burst  ;
	input  [3:0]    Init8_Ar_Cache  ;
	input  [7:0]    Init8_Ar_Id     ;
	input  [7:0]    Init8_Ar_Len    ;
	input  [1:0]    Init8_Ar_Lock   ;
	input  [2:0]    Init8_Ar_Prot   ;
	input  [3:0]    Init8_Ar_Qos    ;
	output          Init8_Ar_Ready  ;
	input  [2:0]    Init8_Ar_Size   ;
	input  [7:0]    Init8_Ar_User   ;
	input           Init8_Ar_Valid  ;
	input  [52:0]   Init8_Aw_Addr   ;
	input  [1:0]    Init8_Aw_Burst  ;
	input  [3:0]    Init8_Aw_Cache  ;
	input  [7:0]    Init8_Aw_Id     ;
	input  [7:0]    Init8_Aw_Len    ;
	input  [1:0]    Init8_Aw_Lock   ;
	input  [2:0]    Init8_Aw_Prot   ;
	input  [3:0]    Init8_Aw_Qos    ;
	output          Init8_Aw_Ready  ;
	input  [2:0]    Init8_Aw_Size   ;
	input  [7:0]    Init8_Aw_User   ;
	input           Init8_Aw_Valid  ;
	output [7:0]    Init8_B_Id      ;
	input           Init8_B_Ready   ;
	output [1:0]    Init8_B_Resp    ;
	output [7:0]    Init8_B_User    ;
	output          Init8_B_Valid   ;
	output [1023:0] Init8_R_Data    ;
	output [7:0]    Init8_R_Id      ;
	output          Init8_R_Last    ;
	input           Init8_R_Ready   ;
	output [1:0]    Init8_R_Resp    ;
	output [7:0]    Init8_R_User    ;
	output          Init8_R_Valid   ;
	input  [1023:0] Init8_W_Data    ;
	input  [7:0]    Init8_W_Id      ;
	input           Init8_W_Last    ;
	output          Init8_W_Ready   ;
	input  [127:0]  Init8_W_Strb    ;
	input           Init8_W_Valid   ;
	input  [52:0]   Init9_Ar_Addr   ;
	input  [1:0]    Init9_Ar_Burst  ;
	input  [3:0]    Init9_Ar_Cache  ;
	input  [7:0]    Init9_Ar_Id     ;
	input  [7:0]    Init9_Ar_Len    ;
	input  [1:0]    Init9_Ar_Lock   ;
	input  [2:0]    Init9_Ar_Prot   ;
	input  [3:0]    Init9_Ar_Qos    ;
	output          Init9_Ar_Ready  ;
	input  [2:0]    Init9_Ar_Size   ;
	input  [7:0]    Init9_Ar_User   ;
	input           Init9_Ar_Valid  ;
	input  [52:0]   Init9_Aw_Addr   ;
	input  [1:0]    Init9_Aw_Burst  ;
	input  [3:0]    Init9_Aw_Cache  ;
	input  [7:0]    Init9_Aw_Id     ;
	input  [7:0]    Init9_Aw_Len    ;
	input  [1:0]    Init9_Aw_Lock   ;
	input  [2:0]    Init9_Aw_Prot   ;
	input  [3:0]    Init9_Aw_Qos    ;
	output          Init9_Aw_Ready  ;
	input  [2:0]    Init9_Aw_Size   ;
	input  [7:0]    Init9_Aw_User   ;
	input           Init9_Aw_Valid  ;
	output [7:0]    Init9_B_Id      ;
	input           Init9_B_Ready   ;
	output [1:0]    Init9_B_Resp    ;
	output [7:0]    Init9_B_User    ;
	output          Init9_B_Valid   ;
	output [1023:0] Init9_R_Data    ;
	output [7:0]    Init9_R_Id      ;
	output          Init9_R_Last    ;
	input           Init9_R_Ready   ;
	output [1:0]    Init9_R_Resp    ;
	output [7:0]    Init9_R_User    ;
	output          Init9_R_Valid   ;
	input  [1023:0] Init9_W_Data    ;
	input  [7:0]    Init9_W_Id      ;
	input           Init9_W_Last    ;
	output          Init9_W_Ready   ;
	input  [127:0]  Init9_W_Strb    ;
	input           Init9_W_Valid   ;
	output [52:0]   Targ0_Ar_Addr   ;
	output [1:0]    Targ0_Ar_Burst  ;
	output [3:0]    Targ0_Ar_Cache  ;
	output [7:0]    Targ0_Ar_Id     ;
	output [7:0]    Targ0_Ar_Len    ;
	output [1:0]    Targ0_Ar_Lock   ;
	output [2:0]    Targ0_Ar_Prot   ;
	output [3:0]    Targ0_Ar_Qos    ;
	input           Targ0_Ar_Ready  ;
	output [2:0]    Targ0_Ar_Size   ;
	output [7:0]    Targ0_Ar_User   ;
	output          Targ0_Ar_Valid  ;
	output [52:0]   Targ0_Aw_Addr   ;
	output [1:0]    Targ0_Aw_Burst  ;
	output [3:0]    Targ0_Aw_Cache  ;
	output [7:0]    Targ0_Aw_Id     ;
	output [7:0]    Targ0_Aw_Len    ;
	output [1:0]    Targ0_Aw_Lock   ;
	output [2:0]    Targ0_Aw_Prot   ;
	output [3:0]    Targ0_Aw_Qos    ;
	input           Targ0_Aw_Ready  ;
	output [2:0]    Targ0_Aw_Size   ;
	output [7:0]    Targ0_Aw_User   ;
	output          Targ0_Aw_Valid  ;
	input  [7:0]    Targ0_B_Id      ;
	output          Targ0_B_Ready   ;
	input  [1:0]    Targ0_B_Resp    ;
	input  [7:0]    Targ0_B_User    ;
	input           Targ0_B_Valid   ;
	input  [1023:0] Targ0_R_Data    ;
	input  [7:0]    Targ0_R_Id      ;
	input           Targ0_R_Last    ;
	output          Targ0_R_Ready   ;
	input  [1:0]    Targ0_R_Resp    ;
	input  [7:0]    Targ0_R_User    ;
	input           Targ0_R_Valid   ;
	output [1023:0] Targ0_W_Data    ;
	output [7:0]    Targ0_W_Id      ;
	output          Targ0_W_Last    ;
	input           Targ0_W_Ready   ;
	output [127:0]  Targ0_W_Strb    ;
	output          Targ0_W_Valid   ;
	output [52:0]   Targ1_Ar_Addr   ;
	output [1:0]    Targ1_Ar_Burst  ;
	output [3:0]    Targ1_Ar_Cache  ;
	output [7:0]    Targ1_Ar_Id     ;
	output [7:0]    Targ1_Ar_Len    ;
	output [1:0]    Targ1_Ar_Lock   ;
	output [2:0]    Targ1_Ar_Prot   ;
	output [3:0]    Targ1_Ar_Qos    ;
	input           Targ1_Ar_Ready  ;
	output [2:0]    Targ1_Ar_Size   ;
	output [7:0]    Targ1_Ar_User   ;
	output          Targ1_Ar_Valid  ;
	output [52:0]   Targ1_Aw_Addr   ;
	output [1:0]    Targ1_Aw_Burst  ;
	output [3:0]    Targ1_Aw_Cache  ;
	output [7:0]    Targ1_Aw_Id     ;
	output [7:0]    Targ1_Aw_Len    ;
	output [1:0]    Targ1_Aw_Lock   ;
	output [2:0]    Targ1_Aw_Prot   ;
	output [3:0]    Targ1_Aw_Qos    ;
	input           Targ1_Aw_Ready  ;
	output [2:0]    Targ1_Aw_Size   ;
	output [7:0]    Targ1_Aw_User   ;
	output          Targ1_Aw_Valid  ;
	input  [7:0]    Targ1_B_Id      ;
	output          Targ1_B_Ready   ;
	input  [1:0]    Targ1_B_Resp    ;
	input  [7:0]    Targ1_B_User    ;
	input           Targ1_B_Valid   ;
	input  [1023:0] Targ1_R_Data    ;
	input  [7:0]    Targ1_R_Id      ;
	input           Targ1_R_Last    ;
	output          Targ1_R_Ready   ;
	input  [1:0]    Targ1_R_Resp    ;
	input  [7:0]    Targ1_R_User    ;
	input           Targ1_R_Valid   ;
	output [1023:0] Targ1_W_Data    ;
	output [7:0]    Targ1_W_Id      ;
	output          Targ1_W_Last    ;
	input           Targ1_W_Ready   ;
	output [127:0]  Targ1_W_Strb    ;
	output          Targ1_W_Valid   ;
	output [52:0]   Targ10_Ar_Addr  ;
	output [1:0]    Targ10_Ar_Burst ;
	output [3:0]    Targ10_Ar_Cache ;
	output [7:0]    Targ10_Ar_Id    ;
	output [7:0]    Targ10_Ar_Len   ;
	output [1:0]    Targ10_Ar_Lock  ;
	output [2:0]    Targ10_Ar_Prot  ;
	output [3:0]    Targ10_Ar_Qos   ;
	input           Targ10_Ar_Ready ;
	output [2:0]    Targ10_Ar_Size  ;
	output [7:0]    Targ10_Ar_User  ;
	output          Targ10_Ar_Valid ;
	output [52:0]   Targ10_Aw_Addr  ;
	output [1:0]    Targ10_Aw_Burst ;
	output [3:0]    Targ10_Aw_Cache ;
	output [7:0]    Targ10_Aw_Id    ;
	output [7:0]    Targ10_Aw_Len   ;
	output [1:0]    Targ10_Aw_Lock  ;
	output [2:0]    Targ10_Aw_Prot  ;
	output [3:0]    Targ10_Aw_Qos   ;
	input           Targ10_Aw_Ready ;
	output [2:0]    Targ10_Aw_Size  ;
	output [7:0]    Targ10_Aw_User  ;
	output          Targ10_Aw_Valid ;
	input  [7:0]    Targ10_B_Id     ;
	output          Targ10_B_Ready  ;
	input  [1:0]    Targ10_B_Resp   ;
	input  [7:0]    Targ10_B_User   ;
	input           Targ10_B_Valid  ;
	input  [1023:0] Targ10_R_Data   ;
	input  [7:0]    Targ10_R_Id     ;
	input           Targ10_R_Last   ;
	output          Targ10_R_Ready  ;
	input  [1:0]    Targ10_R_Resp   ;
	input  [7:0]    Targ10_R_User   ;
	input           Targ10_R_Valid  ;
	output [1023:0] Targ10_W_Data   ;
	output [7:0]    Targ10_W_Id     ;
	output          Targ10_W_Last   ;
	input           Targ10_W_Ready  ;
	output [127:0]  Targ10_W_Strb   ;
	output          Targ10_W_Valid  ;
	output [52:0]   Targ11_Ar_Addr  ;
	output [1:0]    Targ11_Ar_Burst ;
	output [3:0]    Targ11_Ar_Cache ;
	output [7:0]    Targ11_Ar_Id    ;
	output [7:0]    Targ11_Ar_Len   ;
	output [1:0]    Targ11_Ar_Lock  ;
	output [2:0]    Targ11_Ar_Prot  ;
	output [3:0]    Targ11_Ar_Qos   ;
	input           Targ11_Ar_Ready ;
	output [2:0]    Targ11_Ar_Size  ;
	output [7:0]    Targ11_Ar_User  ;
	output          Targ11_Ar_Valid ;
	output [52:0]   Targ11_Aw_Addr  ;
	output [1:0]    Targ11_Aw_Burst ;
	output [3:0]    Targ11_Aw_Cache ;
	output [7:0]    Targ11_Aw_Id    ;
	output [7:0]    Targ11_Aw_Len   ;
	output [1:0]    Targ11_Aw_Lock  ;
	output [2:0]    Targ11_Aw_Prot  ;
	output [3:0]    Targ11_Aw_Qos   ;
	input           Targ11_Aw_Ready ;
	output [2:0]    Targ11_Aw_Size  ;
	output [7:0]    Targ11_Aw_User  ;
	output          Targ11_Aw_Valid ;
	input  [7:0]    Targ11_B_Id     ;
	output          Targ11_B_Ready  ;
	input  [1:0]    Targ11_B_Resp   ;
	input  [7:0]    Targ11_B_User   ;
	input           Targ11_B_Valid  ;
	input  [1023:0] Targ11_R_Data   ;
	input  [7:0]    Targ11_R_Id     ;
	input           Targ11_R_Last   ;
	output          Targ11_R_Ready  ;
	input  [1:0]    Targ11_R_Resp   ;
	input  [7:0]    Targ11_R_User   ;
	input           Targ11_R_Valid  ;
	output [1023:0] Targ11_W_Data   ;
	output [7:0]    Targ11_W_Id     ;
	output          Targ11_W_Last   ;
	input           Targ11_W_Ready  ;
	output [127:0]  Targ11_W_Strb   ;
	output          Targ11_W_Valid  ;
	output [52:0]   Targ2_Ar_Addr   ;
	output [1:0]    Targ2_Ar_Burst  ;
	output [3:0]    Targ2_Ar_Cache  ;
	output [7:0]    Targ2_Ar_Id     ;
	output [7:0]    Targ2_Ar_Len    ;
	output [1:0]    Targ2_Ar_Lock   ;
	output [2:0]    Targ2_Ar_Prot   ;
	output [3:0]    Targ2_Ar_Qos    ;
	input           Targ2_Ar_Ready  ;
	output [2:0]    Targ2_Ar_Size   ;
	output [7:0]    Targ2_Ar_User   ;
	output          Targ2_Ar_Valid  ;
	output [52:0]   Targ2_Aw_Addr   ;
	output [1:0]    Targ2_Aw_Burst  ;
	output [3:0]    Targ2_Aw_Cache  ;
	output [7:0]    Targ2_Aw_Id     ;
	output [7:0]    Targ2_Aw_Len    ;
	output [1:0]    Targ2_Aw_Lock   ;
	output [2:0]    Targ2_Aw_Prot   ;
	output [3:0]    Targ2_Aw_Qos    ;
	input           Targ2_Aw_Ready  ;
	output [2:0]    Targ2_Aw_Size   ;
	output [7:0]    Targ2_Aw_User   ;
	output          Targ2_Aw_Valid  ;
	input  [7:0]    Targ2_B_Id      ;
	output          Targ2_B_Ready   ;
	input  [1:0]    Targ2_B_Resp    ;
	input  [7:0]    Targ2_B_User    ;
	input           Targ2_B_Valid   ;
	input  [1023:0] Targ2_R_Data    ;
	input  [7:0]    Targ2_R_Id      ;
	input           Targ2_R_Last    ;
	output          Targ2_R_Ready   ;
	input  [1:0]    Targ2_R_Resp    ;
	input  [7:0]    Targ2_R_User    ;
	input           Targ2_R_Valid   ;
	output [1023:0] Targ2_W_Data    ;
	output [7:0]    Targ2_W_Id      ;
	output          Targ2_W_Last    ;
	input           Targ2_W_Ready   ;
	output [127:0]  Targ2_W_Strb    ;
	output          Targ2_W_Valid   ;
	output [52:0]   Targ3_Ar_Addr   ;
	output [1:0]    Targ3_Ar_Burst  ;
	output [3:0]    Targ3_Ar_Cache  ;
	output [7:0]    Targ3_Ar_Id     ;
	output [7:0]    Targ3_Ar_Len    ;
	output [1:0]    Targ3_Ar_Lock   ;
	output [2:0]    Targ3_Ar_Prot   ;
	output [3:0]    Targ3_Ar_Qos    ;
	input           Targ3_Ar_Ready  ;
	output [2:0]    Targ3_Ar_Size   ;
	output [7:0]    Targ3_Ar_User   ;
	output          Targ3_Ar_Valid  ;
	output [52:0]   Targ3_Aw_Addr   ;
	output [1:0]    Targ3_Aw_Burst  ;
	output [3:0]    Targ3_Aw_Cache  ;
	output [7:0]    Targ3_Aw_Id     ;
	output [7:0]    Targ3_Aw_Len    ;
	output [1:0]    Targ3_Aw_Lock   ;
	output [2:0]    Targ3_Aw_Prot   ;
	output [3:0]    Targ3_Aw_Qos    ;
	input           Targ3_Aw_Ready  ;
	output [2:0]    Targ3_Aw_Size   ;
	output [7:0]    Targ3_Aw_User   ;
	output          Targ3_Aw_Valid  ;
	input  [7:0]    Targ3_B_Id      ;
	output          Targ3_B_Ready   ;
	input  [1:0]    Targ3_B_Resp    ;
	input  [7:0]    Targ3_B_User    ;
	input           Targ3_B_Valid   ;
	input  [1023:0] Targ3_R_Data    ;
	input  [7:0]    Targ3_R_Id      ;
	input           Targ3_R_Last    ;
	output          Targ3_R_Ready   ;
	input  [1:0]    Targ3_R_Resp    ;
	input  [7:0]    Targ3_R_User    ;
	input           Targ3_R_Valid   ;
	output [1023:0] Targ3_W_Data    ;
	output [7:0]    Targ3_W_Id      ;
	output          Targ3_W_Last    ;
	input           Targ3_W_Ready   ;
	output [127:0]  Targ3_W_Strb    ;
	output          Targ3_W_Valid   ;
	output [52:0]   Targ4_Ar_Addr   ;
	output [1:0]    Targ4_Ar_Burst  ;
	output [3:0]    Targ4_Ar_Cache  ;
	output [7:0]    Targ4_Ar_Id     ;
	output [7:0]    Targ4_Ar_Len    ;
	output [1:0]    Targ4_Ar_Lock   ;
	output [2:0]    Targ4_Ar_Prot   ;
	output [3:0]    Targ4_Ar_Qos    ;
	input           Targ4_Ar_Ready  ;
	output [2:0]    Targ4_Ar_Size   ;
	output [7:0]    Targ4_Ar_User   ;
	output          Targ4_Ar_Valid  ;
	output [52:0]   Targ4_Aw_Addr   ;
	output [1:0]    Targ4_Aw_Burst  ;
	output [3:0]    Targ4_Aw_Cache  ;
	output [7:0]    Targ4_Aw_Id     ;
	output [7:0]    Targ4_Aw_Len    ;
	output [1:0]    Targ4_Aw_Lock   ;
	output [2:0]    Targ4_Aw_Prot   ;
	output [3:0]    Targ4_Aw_Qos    ;
	input           Targ4_Aw_Ready  ;
	output [2:0]    Targ4_Aw_Size   ;
	output [7:0]    Targ4_Aw_User   ;
	output          Targ4_Aw_Valid  ;
	input  [7:0]    Targ4_B_Id      ;
	output          Targ4_B_Ready   ;
	input  [1:0]    Targ4_B_Resp    ;
	input  [7:0]    Targ4_B_User    ;
	input           Targ4_B_Valid   ;
	input  [1023:0] Targ4_R_Data    ;
	input  [7:0]    Targ4_R_Id      ;
	input           Targ4_R_Last    ;
	output          Targ4_R_Ready   ;
	input  [1:0]    Targ4_R_Resp    ;
	input  [7:0]    Targ4_R_User    ;
	input           Targ4_R_Valid   ;
	output [1023:0] Targ4_W_Data    ;
	output [7:0]    Targ4_W_Id      ;
	output          Targ4_W_Last    ;
	input           Targ4_W_Ready   ;
	output [127:0]  Targ4_W_Strb    ;
	output          Targ4_W_Valid   ;
	output [52:0]   Targ5_Ar_Addr   ;
	output [1:0]    Targ5_Ar_Burst  ;
	output [3:0]    Targ5_Ar_Cache  ;
	output [7:0]    Targ5_Ar_Id     ;
	output [7:0]    Targ5_Ar_Len    ;
	output [1:0]    Targ5_Ar_Lock   ;
	output [2:0]    Targ5_Ar_Prot   ;
	output [3:0]    Targ5_Ar_Qos    ;
	input           Targ5_Ar_Ready  ;
	output [2:0]    Targ5_Ar_Size   ;
	output [7:0]    Targ5_Ar_User   ;
	output          Targ5_Ar_Valid  ;
	output [52:0]   Targ5_Aw_Addr   ;
	output [1:0]    Targ5_Aw_Burst  ;
	output [3:0]    Targ5_Aw_Cache  ;
	output [7:0]    Targ5_Aw_Id     ;
	output [7:0]    Targ5_Aw_Len    ;
	output [1:0]    Targ5_Aw_Lock   ;
	output [2:0]    Targ5_Aw_Prot   ;
	output [3:0]    Targ5_Aw_Qos    ;
	input           Targ5_Aw_Ready  ;
	output [2:0]    Targ5_Aw_Size   ;
	output [7:0]    Targ5_Aw_User   ;
	output          Targ5_Aw_Valid  ;
	input  [7:0]    Targ5_B_Id      ;
	output          Targ5_B_Ready   ;
	input  [1:0]    Targ5_B_Resp    ;
	input  [7:0]    Targ5_B_User    ;
	input           Targ5_B_Valid   ;
	input  [1023:0] Targ5_R_Data    ;
	input  [7:0]    Targ5_R_Id      ;
	input           Targ5_R_Last    ;
	output          Targ5_R_Ready   ;
	input  [1:0]    Targ5_R_Resp    ;
	input  [7:0]    Targ5_R_User    ;
	input           Targ5_R_Valid   ;
	output [1023:0] Targ5_W_Data    ;
	output [7:0]    Targ5_W_Id      ;
	output          Targ5_W_Last    ;
	input           Targ5_W_Ready   ;
	output [127:0]  Targ5_W_Strb    ;
	output          Targ5_W_Valid   ;
	output [52:0]   Targ6_Ar_Addr   ;
	output [1:0]    Targ6_Ar_Burst  ;
	output [3:0]    Targ6_Ar_Cache  ;
	output [7:0]    Targ6_Ar_Id     ;
	output [7:0]    Targ6_Ar_Len    ;
	output [1:0]    Targ6_Ar_Lock   ;
	output [2:0]    Targ6_Ar_Prot   ;
	output [3:0]    Targ6_Ar_Qos    ;
	input           Targ6_Ar_Ready  ;
	output [2:0]    Targ6_Ar_Size   ;
	output [7:0]    Targ6_Ar_User   ;
	output          Targ6_Ar_Valid  ;
	output [52:0]   Targ6_Aw_Addr   ;
	output [1:0]    Targ6_Aw_Burst  ;
	output [3:0]    Targ6_Aw_Cache  ;
	output [7:0]    Targ6_Aw_Id     ;
	output [7:0]    Targ6_Aw_Len    ;
	output [1:0]    Targ6_Aw_Lock   ;
	output [2:0]    Targ6_Aw_Prot   ;
	output [3:0]    Targ6_Aw_Qos    ;
	input           Targ6_Aw_Ready  ;
	output [2:0]    Targ6_Aw_Size   ;
	output [7:0]    Targ6_Aw_User   ;
	output          Targ6_Aw_Valid  ;
	input  [7:0]    Targ6_B_Id      ;
	output          Targ6_B_Ready   ;
	input  [1:0]    Targ6_B_Resp    ;
	input  [7:0]    Targ6_B_User    ;
	input           Targ6_B_Valid   ;
	input  [1023:0] Targ6_R_Data    ;
	input  [7:0]    Targ6_R_Id      ;
	input           Targ6_R_Last    ;
	output          Targ6_R_Ready   ;
	input  [1:0]    Targ6_R_Resp    ;
	input  [7:0]    Targ6_R_User    ;
	input           Targ6_R_Valid   ;
	output [1023:0] Targ6_W_Data    ;
	output [7:0]    Targ6_W_Id      ;
	output          Targ6_W_Last    ;
	input           Targ6_W_Ready   ;
	output [127:0]  Targ6_W_Strb    ;
	output          Targ6_W_Valid   ;
	output [52:0]   Targ7_Ar_Addr   ;
	output [1:0]    Targ7_Ar_Burst  ;
	output [3:0]    Targ7_Ar_Cache  ;
	output [7:0]    Targ7_Ar_Id     ;
	output [7:0]    Targ7_Ar_Len    ;
	output [1:0]    Targ7_Ar_Lock   ;
	output [2:0]    Targ7_Ar_Prot   ;
	output [3:0]    Targ7_Ar_Qos    ;
	input           Targ7_Ar_Ready  ;
	output [2:0]    Targ7_Ar_Size   ;
	output [7:0]    Targ7_Ar_User   ;
	output          Targ7_Ar_Valid  ;
	output [52:0]   Targ7_Aw_Addr   ;
	output [1:0]    Targ7_Aw_Burst  ;
	output [3:0]    Targ7_Aw_Cache  ;
	output [7:0]    Targ7_Aw_Id     ;
	output [7:0]    Targ7_Aw_Len    ;
	output [1:0]    Targ7_Aw_Lock   ;
	output [2:0]    Targ7_Aw_Prot   ;
	output [3:0]    Targ7_Aw_Qos    ;
	input           Targ7_Aw_Ready  ;
	output [2:0]    Targ7_Aw_Size   ;
	output [7:0]    Targ7_Aw_User   ;
	output          Targ7_Aw_Valid  ;
	input  [7:0]    Targ7_B_Id      ;
	output          Targ7_B_Ready   ;
	input  [1:0]    Targ7_B_Resp    ;
	input  [7:0]    Targ7_B_User    ;
	input           Targ7_B_Valid   ;
	input  [1023:0] Targ7_R_Data    ;
	input  [7:0]    Targ7_R_Id      ;
	input           Targ7_R_Last    ;
	output          Targ7_R_Ready   ;
	input  [1:0]    Targ7_R_Resp    ;
	input  [7:0]    Targ7_R_User    ;
	input           Targ7_R_Valid   ;
	output [1023:0] Targ7_W_Data    ;
	output [7:0]    Targ7_W_Id      ;
	output          Targ7_W_Last    ;
	input           Targ7_W_Ready   ;
	output [127:0]  Targ7_W_Strb    ;
	output          Targ7_W_Valid   ;
	output [52:0]   Targ8_Ar_Addr   ;
	output [1:0]    Targ8_Ar_Burst  ;
	output [3:0]    Targ8_Ar_Cache  ;
	output [7:0]    Targ8_Ar_Id     ;
	output [7:0]    Targ8_Ar_Len    ;
	output [1:0]    Targ8_Ar_Lock   ;
	output [2:0]    Targ8_Ar_Prot   ;
	output [3:0]    Targ8_Ar_Qos    ;
	input           Targ8_Ar_Ready  ;
	output [2:0]    Targ8_Ar_Size   ;
	output [7:0]    Targ8_Ar_User   ;
	output          Targ8_Ar_Valid  ;
	output [52:0]   Targ8_Aw_Addr   ;
	output [1:0]    Targ8_Aw_Burst  ;
	output [3:0]    Targ8_Aw_Cache  ;
	output [7:0]    Targ8_Aw_Id     ;
	output [7:0]    Targ8_Aw_Len    ;
	output [1:0]    Targ8_Aw_Lock   ;
	output [2:0]    Targ8_Aw_Prot   ;
	output [3:0]    Targ8_Aw_Qos    ;
	input           Targ8_Aw_Ready  ;
	output [2:0]    Targ8_Aw_Size   ;
	output [7:0]    Targ8_Aw_User   ;
	output          Targ8_Aw_Valid  ;
	input  [7:0]    Targ8_B_Id      ;
	output          Targ8_B_Ready   ;
	input  [1:0]    Targ8_B_Resp    ;
	input  [7:0]    Targ8_B_User    ;
	input           Targ8_B_Valid   ;
	input  [1023:0] Targ8_R_Data    ;
	input  [7:0]    Targ8_R_Id      ;
	input           Targ8_R_Last    ;
	output          Targ8_R_Ready   ;
	input  [1:0]    Targ8_R_Resp    ;
	input  [7:0]    Targ8_R_User    ;
	input           Targ8_R_Valid   ;
	output [1023:0] Targ8_W_Data    ;
	output [7:0]    Targ8_W_Id      ;
	output          Targ8_W_Last    ;
	input           Targ8_W_Ready   ;
	output [127:0]  Targ8_W_Strb    ;
	output          Targ8_W_Valid   ;
	output [52:0]   Targ9_Ar_Addr   ;
	output [1:0]    Targ9_Ar_Burst  ;
	output [3:0]    Targ9_Ar_Cache  ;
	output [7:0]    Targ9_Ar_Id     ;
	output [7:0]    Targ9_Ar_Len    ;
	output [1:0]    Targ9_Ar_Lock   ;
	output [2:0]    Targ9_Ar_Prot   ;
	output [3:0]    Targ9_Ar_Qos    ;
	input           Targ9_Ar_Ready  ;
	output [2:0]    Targ9_Ar_Size   ;
	output [7:0]    Targ9_Ar_User   ;
	output          Targ9_Ar_Valid  ;
	output [52:0]   Targ9_Aw_Addr   ;
	output [1:0]    Targ9_Aw_Burst  ;
	output [3:0]    Targ9_Aw_Cache  ;
	output [7:0]    Targ9_Aw_Id     ;
	output [7:0]    Targ9_Aw_Len    ;
	output [1:0]    Targ9_Aw_Lock   ;
	output [2:0]    Targ9_Aw_Prot   ;
	output [3:0]    Targ9_Aw_Qos    ;
	input           Targ9_Aw_Ready  ;
	output [2:0]    Targ9_Aw_Size   ;
	output [7:0]    Targ9_Aw_User   ;
	output          Targ9_Aw_Valid  ;
	input  [7:0]    Targ9_B_Id      ;
	output          Targ9_B_Ready   ;
	input  [1:0]    Targ9_B_Resp    ;
	input  [7:0]    Targ9_B_User    ;
	input           Targ9_B_Valid   ;
	input  [1023:0] Targ9_R_Data    ;
	input  [7:0]    Targ9_R_Id      ;
	input           Targ9_R_Last    ;
	output          Targ9_R_Ready   ;
	input  [1:0]    Targ9_R_Resp    ;
	input  [7:0]    Targ9_R_User    ;
	input           Targ9_R_Valid   ;
	output [1023:0] Targ9_W_Data    ;
	output [7:0]    Targ9_W_Id      ;
	output          Targ9_W_Last    ;
	input           Targ9_W_Ready   ;
	output [127:0]  Targ9_W_Strb    ;
	output          Targ9_W_Valid   ;
	input           noc_arstn       ;
	input           node0_aclk      ;
	input           node10_aclk     ;
	input           node11_aclk     ;
	input           node1_aclk      ;
	input           node2_aclk      ;
	input           node3_aclk      ;
	input           node4_aclk      ;
	input           node5_aclk      ;
	input           node6_aclk      ;
	input           node7_aclk      ;
	input           node8_aclk      ;
	input           node9_aclk      ;
	input           tm              ;
endmodule



        
/* verilator lint_off WIDTH */        
module newComponent 
   (
   AXI_4_53_1024_8_withQOS_noREGION.inward Init11,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init7,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init6,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init5,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init4,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init3,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init2,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init1,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init0,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init9,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init8,
   AXI_4_53_1024_8_withQOS_noREGION.inward Init10,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ9,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ8,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ5,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ4,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ7,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ6,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ1,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ0,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ3,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ2,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ11,
   AXI_4_53_1024_8_withQOS_noREGION.outward Targ10
   );

   logic  unbound;


    Specification_Architecture_Structure verilognewComponent
      (
        .Init11_Ar_Addr(Init11.ARADDR),
        .Init11_W_Ready(Init11.WREADY),
        .Init11_Aw_Valid(Init11.AWVALID),
        .Init11_Ar_Qos(Init11.ARQOS),
        .Init11_Ar_Id(Init11.ARID),
        .Init11_R_User(Init11.RUSER),
        .Init11_Aw_Lock(Init11.AWLOCK),
        .Init11_Ar_Lock(Init11.ARLOCK),
        .Init11_Aw_Id(Init11.AWID),
        .Init11_Ar_Len(Init11.ARLEN),
        .Init11_Ar_User(Init11.ARUSER),
        .Init11_B_Id(Init11.BID),
        .Init11_W_Valid(Init11.WVALID),
        .Init11_B_Ready(Init11.BREADY),
        .Init11_W_Data(Init11.WDATA),
        .Init11_R_Valid(Init11.RVALID),
        .Init11_R_Data(Init11.RDATA),
        .Init11_R_Id(Init11.RID),
        .Init11_B_Resp(Init11.BRESP),
        .Init11_Aw_Size(Init11.AWSIZE),
        .Init11_Aw_Addr(Init11.AWADDR),
        .Init11_Aw_Cache(Init11.AWCACHE),
        .Init11_W_Last(Init11.WLAST),
        .Init11_R_Ready(Init11.RREADY),
        .Init11_Ar_Ready(Init11.ARREADY),
        .Init11_Ar_Cache(Init11.ARCACHE),
        .Init11_R_Last(Init11.RLAST),
        .Init11_Aw_Qos(Init11.AWQOS),
        .Init11_Ar_Valid(Init11.ARVALID),
        .Init11_Aw_User(Init11.AWUSER),
        .Init11_Ar_Size(Init11.ARSIZE),
        .Init11_Aw_Ready(Init11.AWREADY),
        .Init11_W_Id(Init11.WID),
        .Init11_B_User(Init11.BUSER),
        .Init11_Ar_Prot(Init11.ARPROT),
        .Init11_Ar_Burst(Init11.ARBURST),
        .Init11_R_Resp(Init11.RRESP),
        .Init11_Aw_Len(Init11.AWLEN),
        .Init11_Aw_Prot(Init11.AWPROT),
        .Init11_W_Strb(Init11.WSTRB),
        .Init11_Aw_Burst(Init11.AWBURST),
        .Init11_B_Valid(Init11.BVALID),
        .node11_aclk(Targ11.ACLK),
        .noc_arstn(Targ10.ARESETn),
        .Init7_Ar_Addr(Init7.ARADDR),
        .Init7_W_Ready(Init7.WREADY),
        .Init7_Aw_Valid(Init7.AWVALID),
        .Init7_Ar_Qos(Init7.ARQOS),
        .Init7_Ar_Id(Init7.ARID),
        .Init7_R_User(Init7.RUSER),
        .Init7_Aw_Lock(Init7.AWLOCK),
        .Init7_Ar_Lock(Init7.ARLOCK),
        .Init7_Aw_Id(Init7.AWID),
        .Init7_Ar_Len(Init7.ARLEN),
        .Init7_Ar_User(Init7.ARUSER),
        .Init7_B_Id(Init7.BID),
        .Init7_W_Valid(Init7.WVALID),
        .Init7_B_Ready(Init7.BREADY),
        .Init7_W_Data(Init7.WDATA),
        .Init7_R_Valid(Init7.RVALID),
        .Init7_R_Data(Init7.RDATA),
        .Init7_R_Id(Init7.RID),
        .Init7_B_Resp(Init7.BRESP),
        .Init7_Aw_Size(Init7.AWSIZE),
        .Init7_Aw_Addr(Init7.AWADDR),
        .Init7_Aw_Cache(Init7.AWCACHE),
        .Init7_W_Last(Init7.WLAST),
        .Init7_R_Ready(Init7.RREADY),
        .Init7_Ar_Ready(Init7.ARREADY),
        .Init7_Ar_Cache(Init7.ARCACHE),
        .Init7_R_Last(Init7.RLAST),
        .Init7_Aw_Qos(Init7.AWQOS),
        .Init7_Ar_Valid(Init7.ARVALID),
        .Init7_Aw_User(Init7.AWUSER),
        .Init7_Ar_Size(Init7.ARSIZE),
        .Init7_Aw_Ready(Init7.AWREADY),
        .Init7_W_Id(Init7.WID),
        .Init7_B_User(Init7.BUSER),
        .Init7_Ar_Prot(Init7.ARPROT),
        .Init7_Ar_Burst(Init7.ARBURST),
        .Init7_R_Resp(Init7.RRESP),
        .Init7_Aw_Len(Init7.AWLEN),
        .Init7_Aw_Prot(Init7.AWPROT),
        .Init7_W_Strb(Init7.WSTRB),
        .Init7_Aw_Burst(Init7.AWBURST),
        .Init7_B_Valid(Init7.BVALID),
        .node7_aclk(Targ7.ACLK),
        .Init6_Ar_Addr(Init6.ARADDR),
        .Init6_W_Ready(Init6.WREADY),
        .Init6_Aw_Valid(Init6.AWVALID),
        .Init6_Ar_Qos(Init6.ARQOS),
        .Init6_Ar_Id(Init6.ARID),
        .Init6_R_User(Init6.RUSER),
        .Init6_Aw_Lock(Init6.AWLOCK),
        .Init6_Ar_Lock(Init6.ARLOCK),
        .Init6_Aw_Id(Init6.AWID),
        .Init6_Ar_Len(Init6.ARLEN),
        .Init6_Ar_User(Init6.ARUSER),
        .Init6_B_Id(Init6.BID),
        .Init6_W_Valid(Init6.WVALID),
        .Init6_B_Ready(Init6.BREADY),
        .Init6_W_Data(Init6.WDATA),
        .Init6_R_Valid(Init6.RVALID),
        .Init6_R_Data(Init6.RDATA),
        .Init6_R_Id(Init6.RID),
        .Init6_B_Resp(Init6.BRESP),
        .Init6_Aw_Size(Init6.AWSIZE),
        .Init6_Aw_Addr(Init6.AWADDR),
        .Init6_Aw_Cache(Init6.AWCACHE),
        .Init6_W_Last(Init6.WLAST),
        .Init6_R_Ready(Init6.RREADY),
        .Init6_Ar_Ready(Init6.ARREADY),
        .Init6_Ar_Cache(Init6.ARCACHE),
        .Init6_R_Last(Init6.RLAST),
        .Init6_Aw_Qos(Init6.AWQOS),
        .Init6_Ar_Valid(Init6.ARVALID),
        .Init6_Aw_User(Init6.AWUSER),
        .Init6_Ar_Size(Init6.ARSIZE),
        .Init6_Aw_Ready(Init6.AWREADY),
        .Init6_W_Id(Init6.WID),
        .Init6_B_User(Init6.BUSER),
        .Init6_Ar_Prot(Init6.ARPROT),
        .Init6_Ar_Burst(Init6.ARBURST),
        .Init6_R_Resp(Init6.RRESP),
        .Init6_Aw_Len(Init6.AWLEN),
        .Init6_Aw_Prot(Init6.AWPROT),
        .Init6_W_Strb(Init6.WSTRB),
        .Init6_Aw_Burst(Init6.AWBURST),
        .Init6_B_Valid(Init6.BVALID),
        .node6_aclk(Targ6.ACLK),
        .Init5_Ar_Addr(Init5.ARADDR),
        .Init5_W_Ready(Init5.WREADY),
        .Init5_Aw_Valid(Init5.AWVALID),
        .Init5_Ar_Qos(Init5.ARQOS),
        .Init5_Ar_Id(Init5.ARID),
        .Init5_R_User(Init5.RUSER),
        .Init5_Aw_Lock(Init5.AWLOCK),
        .Init5_Ar_Lock(Init5.ARLOCK),
        .Init5_Aw_Id(Init5.AWID),
        .Init5_Ar_Len(Init5.ARLEN),
        .Init5_Ar_User(Init5.ARUSER),
        .Init5_B_Id(Init5.BID),
        .Init5_W_Valid(Init5.WVALID),
        .Init5_B_Ready(Init5.BREADY),
        .Init5_W_Data(Init5.WDATA),
        .Init5_R_Valid(Init5.RVALID),
        .Init5_R_Data(Init5.RDATA),
        .Init5_R_Id(Init5.RID),
        .Init5_B_Resp(Init5.BRESP),
        .Init5_Aw_Size(Init5.AWSIZE),
        .Init5_Aw_Addr(Init5.AWADDR),
        .Init5_Aw_Cache(Init5.AWCACHE),
        .Init5_W_Last(Init5.WLAST),
        .Init5_R_Ready(Init5.RREADY),
        .Init5_Ar_Ready(Init5.ARREADY),
        .Init5_Ar_Cache(Init5.ARCACHE),
        .Init5_R_Last(Init5.RLAST),
        .Init5_Aw_Qos(Init5.AWQOS),
        .Init5_Ar_Valid(Init5.ARVALID),
        .Init5_Aw_User(Init5.AWUSER),
        .Init5_Ar_Size(Init5.ARSIZE),
        .Init5_Aw_Ready(Init5.AWREADY),
        .Init5_W_Id(Init5.WID),
        .Init5_B_User(Init5.BUSER),
        .Init5_Ar_Prot(Init5.ARPROT),
        .Init5_Ar_Burst(Init5.ARBURST),
        .Init5_R_Resp(Init5.RRESP),
        .Init5_Aw_Len(Init5.AWLEN),
        .Init5_Aw_Prot(Init5.AWPROT),
        .Init5_W_Strb(Init5.WSTRB),
        .Init5_Aw_Burst(Init5.AWBURST),
        .Init5_B_Valid(Init5.BVALID),
        .node5_aclk(Targ5.ACLK),
        .Init4_Ar_Addr(Init4.ARADDR),
        .Init4_W_Ready(Init4.WREADY),
        .Init4_Aw_Valid(Init4.AWVALID),
        .Init4_Ar_Qos(Init4.ARQOS),
        .Init4_Ar_Id(Init4.ARID),
        .Init4_R_User(Init4.RUSER),
        .Init4_Aw_Lock(Init4.AWLOCK),
        .Init4_Ar_Lock(Init4.ARLOCK),
        .Init4_Aw_Id(Init4.AWID),
        .Init4_Ar_Len(Init4.ARLEN),
        .Init4_Ar_User(Init4.ARUSER),
        .Init4_B_Id(Init4.BID),
        .Init4_W_Valid(Init4.WVALID),
        .Init4_B_Ready(Init4.BREADY),
        .Init4_W_Data(Init4.WDATA),
        .Init4_R_Valid(Init4.RVALID),
        .Init4_R_Data(Init4.RDATA),
        .Init4_R_Id(Init4.RID),
        .Init4_B_Resp(Init4.BRESP),
        .Init4_Aw_Size(Init4.AWSIZE),
        .Init4_Aw_Addr(Init4.AWADDR),
        .Init4_Aw_Cache(Init4.AWCACHE),
        .Init4_W_Last(Init4.WLAST),
        .Init4_R_Ready(Init4.RREADY),
        .Init4_Ar_Ready(Init4.ARREADY),
        .Init4_Ar_Cache(Init4.ARCACHE),
        .Init4_R_Last(Init4.RLAST),
        .Init4_Aw_Qos(Init4.AWQOS),
        .Init4_Ar_Valid(Init4.ARVALID),
        .Init4_Aw_User(Init4.AWUSER),
        .Init4_Ar_Size(Init4.ARSIZE),
        .Init4_Aw_Ready(Init4.AWREADY),
        .Init4_W_Id(Init4.WID),
        .Init4_B_User(Init4.BUSER),
        .Init4_Ar_Prot(Init4.ARPROT),
        .Init4_Ar_Burst(Init4.ARBURST),
        .Init4_R_Resp(Init4.RRESP),
        .Init4_Aw_Len(Init4.AWLEN),
        .Init4_Aw_Prot(Init4.AWPROT),
        .Init4_W_Strb(Init4.WSTRB),
        .Init4_Aw_Burst(Init4.AWBURST),
        .Init4_B_Valid(Init4.BVALID),
        .node4_aclk(Targ4.ACLK),
        .Init3_Ar_Addr(Init3.ARADDR),
        .Init3_W_Ready(Init3.WREADY),
        .Init3_Aw_Valid(Init3.AWVALID),
        .Init3_Ar_Qos(Init3.ARQOS),
        .Init3_Ar_Id(Init3.ARID),
        .Init3_R_User(Init3.RUSER),
        .Init3_Aw_Lock(Init3.AWLOCK),
        .Init3_Ar_Lock(Init3.ARLOCK),
        .Init3_Aw_Id(Init3.AWID),
        .Init3_Ar_Len(Init3.ARLEN),
        .Init3_Ar_User(Init3.ARUSER),
        .Init3_B_Id(Init3.BID),
        .Init3_W_Valid(Init3.WVALID),
        .Init3_B_Ready(Init3.BREADY),
        .Init3_W_Data(Init3.WDATA),
        .Init3_R_Valid(Init3.RVALID),
        .Init3_R_Data(Init3.RDATA),
        .Init3_R_Id(Init3.RID),
        .Init3_B_Resp(Init3.BRESP),
        .Init3_Aw_Size(Init3.AWSIZE),
        .Init3_Aw_Addr(Init3.AWADDR),
        .Init3_Aw_Cache(Init3.AWCACHE),
        .Init3_W_Last(Init3.WLAST),
        .Init3_R_Ready(Init3.RREADY),
        .Init3_Ar_Ready(Init3.ARREADY),
        .Init3_Ar_Cache(Init3.ARCACHE),
        .Init3_R_Last(Init3.RLAST),
        .Init3_Aw_Qos(Init3.AWQOS),
        .Init3_Ar_Valid(Init3.ARVALID),
        .Init3_Aw_User(Init3.AWUSER),
        .Init3_Ar_Size(Init3.ARSIZE),
        .Init3_Aw_Ready(Init3.AWREADY),
        .Init3_W_Id(Init3.WID),
        .Init3_B_User(Init3.BUSER),
        .Init3_Ar_Prot(Init3.ARPROT),
        .Init3_Ar_Burst(Init3.ARBURST),
        .Init3_R_Resp(Init3.RRESP),
        .Init3_Aw_Len(Init3.AWLEN),
        .Init3_Aw_Prot(Init3.AWPROT),
        .Init3_W_Strb(Init3.WSTRB),
        .Init3_Aw_Burst(Init3.AWBURST),
        .Init3_B_Valid(Init3.BVALID),
        .node3_aclk(Targ3.ACLK),
        .Init2_Ar_Addr(Init2.ARADDR),
        .Init2_W_Ready(Init2.WREADY),
        .Init2_Aw_Valid(Init2.AWVALID),
        .Init2_Ar_Qos(Init2.ARQOS),
        .Init2_Ar_Id(Init2.ARID),
        .Init2_R_User(Init2.RUSER),
        .Init2_Aw_Lock(Init2.AWLOCK),
        .Init2_Ar_Lock(Init2.ARLOCK),
        .Init2_Aw_Id(Init2.AWID),
        .Init2_Ar_Len(Init2.ARLEN),
        .Init2_Ar_User(Init2.ARUSER),
        .Init2_B_Id(Init2.BID),
        .Init2_W_Valid(Init2.WVALID),
        .Init2_B_Ready(Init2.BREADY),
        .Init2_W_Data(Init2.WDATA),
        .Init2_R_Valid(Init2.RVALID),
        .Init2_R_Data(Init2.RDATA),
        .Init2_R_Id(Init2.RID),
        .Init2_B_Resp(Init2.BRESP),
        .Init2_Aw_Size(Init2.AWSIZE),
        .Init2_Aw_Addr(Init2.AWADDR),
        .Init2_Aw_Cache(Init2.AWCACHE),
        .Init2_W_Last(Init2.WLAST),
        .Init2_R_Ready(Init2.RREADY),
        .Init2_Ar_Ready(Init2.ARREADY),
        .Init2_Ar_Cache(Init2.ARCACHE),
        .Init2_R_Last(Init2.RLAST),
        .Init2_Aw_Qos(Init2.AWQOS),
        .Init2_Ar_Valid(Init2.ARVALID),
        .Init2_Aw_User(Init2.AWUSER),
        .Init2_Ar_Size(Init2.ARSIZE),
        .Init2_Aw_Ready(Init2.AWREADY),
        .Init2_W_Id(Init2.WID),
        .Init2_B_User(Init2.BUSER),
        .Init2_Ar_Prot(Init2.ARPROT),
        .Init2_Ar_Burst(Init2.ARBURST),
        .Init2_R_Resp(Init2.RRESP),
        .Init2_Aw_Len(Init2.AWLEN),
        .Init2_Aw_Prot(Init2.AWPROT),
        .Init2_W_Strb(Init2.WSTRB),
        .Init2_Aw_Burst(Init2.AWBURST),
        .Init2_B_Valid(Init2.BVALID),
        .node2_aclk(Targ2.ACLK),
        .Init1_Ar_Addr(Init1.ARADDR),
        .Init1_W_Ready(Init1.WREADY),
        .Init1_Aw_Valid(Init1.AWVALID),
        .Init1_Ar_Qos(Init1.ARQOS),
        .Init1_Ar_Id(Init1.ARID),
        .Init1_R_User(Init1.RUSER),
        .Init1_Aw_Lock(Init1.AWLOCK),
        .Init1_Ar_Lock(Init1.ARLOCK),
        .Init1_Aw_Id(Init1.AWID),
        .Init1_Ar_Len(Init1.ARLEN),
        .Init1_Ar_User(Init1.ARUSER),
        .Init1_B_Id(Init1.BID),
        .Init1_W_Valid(Init1.WVALID),
        .Init1_B_Ready(Init1.BREADY),
        .Init1_W_Data(Init1.WDATA),
        .Init1_R_Valid(Init1.RVALID),
        .Init1_R_Data(Init1.RDATA),
        .Init1_R_Id(Init1.RID),
        .Init1_B_Resp(Init1.BRESP),
        .Init1_Aw_Size(Init1.AWSIZE),
        .Init1_Aw_Addr(Init1.AWADDR),
        .Init1_Aw_Cache(Init1.AWCACHE),
        .Init1_W_Last(Init1.WLAST),
        .Init1_R_Ready(Init1.RREADY),
        .Init1_Ar_Ready(Init1.ARREADY),
        .Init1_Ar_Cache(Init1.ARCACHE),
        .Init1_R_Last(Init1.RLAST),
        .Init1_Aw_Qos(Init1.AWQOS),
        .Init1_Ar_Valid(Init1.ARVALID),
        .Init1_Aw_User(Init1.AWUSER),
        .Init1_Ar_Size(Init1.ARSIZE),
        .Init1_Aw_Ready(Init1.AWREADY),
        .Init1_W_Id(Init1.WID),
        .Init1_B_User(Init1.BUSER),
        .Init1_Ar_Prot(Init1.ARPROT),
        .Init1_Ar_Burst(Init1.ARBURST),
        .Init1_R_Resp(Init1.RRESP),
        .Init1_Aw_Len(Init1.AWLEN),
        .Init1_Aw_Prot(Init1.AWPROT),
        .Init1_W_Strb(Init1.WSTRB),
        .Init1_Aw_Burst(Init1.AWBURST),
        .Init1_B_Valid(Init1.BVALID),
        .node1_aclk(Targ1.ACLK),
        .Init0_Ar_Addr(Init0.ARADDR),
        .Init0_W_Ready(Init0.WREADY),
        .Init0_Aw_Valid(Init0.AWVALID),
        .Init0_Ar_Qos(Init0.ARQOS),
        .Init0_Ar_Id(Init0.ARID),
        .Init0_R_User(Init0.RUSER),
        .Init0_Aw_Lock(Init0.AWLOCK),
        .Init0_Ar_Lock(Init0.ARLOCK),
        .Init0_Aw_Id(Init0.AWID),
        .Init0_Ar_Len(Init0.ARLEN),
        .Init0_Ar_User(Init0.ARUSER),
        .Init0_B_Id(Init0.BID),
        .Init0_W_Valid(Init0.WVALID),
        .Init0_B_Ready(Init0.BREADY),
        .Init0_W_Data(Init0.WDATA),
        .Init0_R_Valid(Init0.RVALID),
        .Init0_R_Data(Init0.RDATA),
        .Init0_R_Id(Init0.RID),
        .Init0_B_Resp(Init0.BRESP),
        .Init0_Aw_Size(Init0.AWSIZE),
        .Init0_Aw_Addr(Init0.AWADDR),
        .Init0_Aw_Cache(Init0.AWCACHE),
        .Init0_W_Last(Init0.WLAST),
        .Init0_R_Ready(Init0.RREADY),
        .Init0_Ar_Ready(Init0.ARREADY),
        .Init0_Ar_Cache(Init0.ARCACHE),
        .Init0_R_Last(Init0.RLAST),
        .Init0_Aw_Qos(Init0.AWQOS),
        .Init0_Ar_Valid(Init0.ARVALID),
        .Init0_Aw_User(Init0.AWUSER),
        .Init0_Ar_Size(Init0.ARSIZE),
        .Init0_Aw_Ready(Init0.AWREADY),
        .Init0_W_Id(Init0.WID),
        .Init0_B_User(Init0.BUSER),
        .Init0_Ar_Prot(Init0.ARPROT),
        .Init0_Ar_Burst(Init0.ARBURST),
        .Init0_R_Resp(Init0.RRESP),
        .Init0_Aw_Len(Init0.AWLEN),
        .Init0_Aw_Prot(Init0.AWPROT),
        .Init0_W_Strb(Init0.WSTRB),
        .Init0_Aw_Burst(Init0.AWBURST),
        .Init0_B_Valid(Init0.BVALID),
        .node0_aclk(Targ0.ACLK),
        .Init9_Ar_Addr(Init9.ARADDR),
        .Init9_W_Ready(Init9.WREADY),
        .Init9_Aw_Valid(Init9.AWVALID),
        .Init9_Ar_Qos(Init9.ARQOS),
        .Init9_Ar_Id(Init9.ARID),
        .Init9_R_User(Init9.RUSER),
        .Init9_Aw_Lock(Init9.AWLOCK),
        .Init9_Ar_Lock(Init9.ARLOCK),
        .Init9_Aw_Id(Init9.AWID),
        .Init9_Ar_Len(Init9.ARLEN),
        .Init9_Ar_User(Init9.ARUSER),
        .Init9_B_Id(Init9.BID),
        .Init9_W_Valid(Init9.WVALID),
        .Init9_B_Ready(Init9.BREADY),
        .Init9_W_Data(Init9.WDATA),
        .Init9_R_Valid(Init9.RVALID),
        .Init9_R_Data(Init9.RDATA),
        .Init9_R_Id(Init9.RID),
        .Init9_B_Resp(Init9.BRESP),
        .Init9_Aw_Size(Init9.AWSIZE),
        .Init9_Aw_Addr(Init9.AWADDR),
        .Init9_Aw_Cache(Init9.AWCACHE),
        .Init9_W_Last(Init9.WLAST),
        .Init9_R_Ready(Init9.RREADY),
        .Init9_Ar_Ready(Init9.ARREADY),
        .Init9_Ar_Cache(Init9.ARCACHE),
        .Init9_R_Last(Init9.RLAST),
        .Init9_Aw_Qos(Init9.AWQOS),
        .Init9_Ar_Valid(Init9.ARVALID),
        .Init9_Aw_User(Init9.AWUSER),
        .Init9_Ar_Size(Init9.ARSIZE),
        .Init9_Aw_Ready(Init9.AWREADY),
        .Init9_W_Id(Init9.WID),
        .Init9_B_User(Init9.BUSER),
        .Init9_Ar_Prot(Init9.ARPROT),
        .Init9_Ar_Burst(Init9.ARBURST),
        .Init9_R_Resp(Init9.RRESP),
        .Init9_Aw_Len(Init9.AWLEN),
        .Init9_Aw_Prot(Init9.AWPROT),
        .Init9_W_Strb(Init9.WSTRB),
        .Init9_Aw_Burst(Init9.AWBURST),
        .Init9_B_Valid(Init9.BVALID),
        .node9_aclk(Targ9.ACLK),
        .Init8_Ar_Addr(Init8.ARADDR),
        .Init8_W_Ready(Init8.WREADY),
        .Init8_Aw_Valid(Init8.AWVALID),
        .Init8_Ar_Qos(Init8.ARQOS),
        .Init8_Ar_Id(Init8.ARID),
        .Init8_R_User(Init8.RUSER),
        .Init8_Aw_Lock(Init8.AWLOCK),
        .Init8_Ar_Lock(Init8.ARLOCK),
        .Init8_Aw_Id(Init8.AWID),
        .Init8_Ar_Len(Init8.ARLEN),
        .Init8_Ar_User(Init8.ARUSER),
        .Init8_B_Id(Init8.BID),
        .Init8_W_Valid(Init8.WVALID),
        .Init8_B_Ready(Init8.BREADY),
        .Init8_W_Data(Init8.WDATA),
        .Init8_R_Valid(Init8.RVALID),
        .Init8_R_Data(Init8.RDATA),
        .Init8_R_Id(Init8.RID),
        .Init8_B_Resp(Init8.BRESP),
        .Init8_Aw_Size(Init8.AWSIZE),
        .Init8_Aw_Addr(Init8.AWADDR),
        .Init8_Aw_Cache(Init8.AWCACHE),
        .Init8_W_Last(Init8.WLAST),
        .Init8_R_Ready(Init8.RREADY),
        .Init8_Ar_Ready(Init8.ARREADY),
        .Init8_Ar_Cache(Init8.ARCACHE),
        .Init8_R_Last(Init8.RLAST),
        .Init8_Aw_Qos(Init8.AWQOS),
        .Init8_Ar_Valid(Init8.ARVALID),
        .Init8_Aw_User(Init8.AWUSER),
        .Init8_Ar_Size(Init8.ARSIZE),
        .Init8_Aw_Ready(Init8.AWREADY),
        .Init8_W_Id(Init8.WID),
        .Init8_B_User(Init8.BUSER),
        .Init8_Ar_Prot(Init8.ARPROT),
        .Init8_Ar_Burst(Init8.ARBURST),
        .Init8_R_Resp(Init8.RRESP),
        .Init8_Aw_Len(Init8.AWLEN),
        .Init8_Aw_Prot(Init8.AWPROT),
        .Init8_W_Strb(Init8.WSTRB),
        .Init8_Aw_Burst(Init8.AWBURST),
        .Init8_B_Valid(Init8.BVALID),
        .node8_aclk(Targ8.ACLK),
        .Init10_Ar_Addr(Init10.ARADDR),
        .Init10_W_Ready(Init10.WREADY),
        .Init10_Aw_Valid(Init10.AWVALID),
        .Init10_Ar_Qos(Init10.ARQOS),
        .Init10_Ar_Id(Init10.ARID),
        .Init10_R_User(Init10.RUSER),
        .Init10_Aw_Lock(Init10.AWLOCK),
        .Init10_Ar_Lock(Init10.ARLOCK),
        .Init10_Aw_Id(Init10.AWID),
        .Init10_Ar_Len(Init10.ARLEN),
        .Init10_Ar_User(Init10.ARUSER),
        .Init10_B_Id(Init10.BID),
        .Init10_W_Valid(Init10.WVALID),
        .Init10_B_Ready(Init10.BREADY),
        .Init10_W_Data(Init10.WDATA),
        .Init10_R_Valid(Init10.RVALID),
        .Init10_R_Data(Init10.RDATA),
        .Init10_R_Id(Init10.RID),
        .Init10_B_Resp(Init10.BRESP),
        .Init10_Aw_Size(Init10.AWSIZE),
        .Init10_Aw_Addr(Init10.AWADDR),
        .Init10_Aw_Cache(Init10.AWCACHE),
        .Init10_W_Last(Init10.WLAST),
        .Init10_R_Ready(Init10.RREADY),
        .Init10_Ar_Ready(Init10.ARREADY),
        .Init10_Ar_Cache(Init10.ARCACHE),
        .Init10_R_Last(Init10.RLAST),
        .Init10_Aw_Qos(Init10.AWQOS),
        .Init10_Ar_Valid(Init10.ARVALID),
        .Init10_Aw_User(Init10.AWUSER),
        .Init10_Ar_Size(Init10.ARSIZE),
        .Init10_Aw_Ready(Init10.AWREADY),
        .Init10_W_Id(Init10.WID),
        .Init10_B_User(Init10.BUSER),
        .Init10_Ar_Prot(Init10.ARPROT),
        .Init10_Ar_Burst(Init10.ARBURST),
        .Init10_R_Resp(Init10.RRESP),
        .Init10_Aw_Len(Init10.AWLEN),
        .Init10_Aw_Prot(Init10.AWPROT),
        .Init10_W_Strb(Init10.WSTRB),
        .Init10_Aw_Burst(Init10.AWBURST),
        .Init10_B_Valid(Init10.BVALID),
        .node10_aclk(Targ10.ACLK),
        .Targ9_Ar_Addr(Targ9.ARADDR),
        .Targ9_W_Ready(Targ9.WREADY),
        .Targ9_Aw_Valid(Targ9.AWVALID),
        .Targ9_Ar_Qos(Targ9.ARQOS),
        .Targ9_Ar_Id(Targ9.ARID),
        .Targ9_R_User(Targ9.RUSER),
        .Targ9_Aw_Lock(Targ9.AWLOCK),
        .Targ9_Ar_Lock(Targ9.ARLOCK),
        .Targ9_Aw_Id(Targ9.AWID),
        .Targ9_Ar_Len(Targ9.ARLEN),
        .Targ9_Ar_User(Targ9.ARUSER),
        .Targ9_B_Id(Targ9.BID),
        .Targ9_W_Valid(Targ9.WVALID),
        .Targ9_B_Ready(Targ9.BREADY),
        .Targ9_W_Data(Targ9.WDATA),
        .Targ9_R_Valid(Targ9.RVALID),
        .Targ9_R_Data(Targ9.RDATA),
        .Targ9_R_Id(Targ9.RID),
        .Targ9_B_Resp(Targ9.BRESP),
        .Targ9_Aw_Size(Targ9.AWSIZE),
        .Targ9_Aw_Addr(Targ9.AWADDR),
        .Targ9_Aw_Cache(Targ9.AWCACHE),
        .Targ9_W_Last(Targ9.WLAST),
        .Targ9_R_Ready(Targ9.RREADY),
        .Targ9_Ar_Ready(Targ9.ARREADY),
        .Targ9_Ar_Cache(Targ9.ARCACHE),
        .Targ9_R_Last(Targ9.RLAST),
        .Targ9_Aw_Qos(Targ9.AWQOS),
        .Targ9_Ar_Valid(Targ9.ARVALID),
        .Targ9_Aw_User(Targ9.AWUSER),
        .Targ9_Ar_Size(Targ9.ARSIZE),
        .Targ9_Aw_Ready(Targ9.AWREADY),
        .Targ9_W_Id(Targ9.WID),
        .Targ9_B_User(Targ9.BUSER),
        .Targ9_Ar_Prot(Targ9.ARPROT),
        .Targ9_Ar_Burst(Targ9.ARBURST),
        .Targ9_R_Resp(Targ9.RRESP),
        .Targ9_Aw_Len(Targ9.AWLEN),
        .Targ9_Aw_Prot(Targ9.AWPROT),
        .Targ9_W_Strb(Targ9.WSTRB),
        .Targ9_Aw_Burst(Targ9.AWBURST),
        .Targ9_B_Valid(Targ9.BVALID),
        .Targ8_Ar_Addr(Targ8.ARADDR),
        .Targ8_W_Ready(Targ8.WREADY),
        .Targ8_Aw_Valid(Targ8.AWVALID),
        .Targ8_Ar_Qos(Targ8.ARQOS),
        .Targ8_Ar_Id(Targ8.ARID),
        .Targ8_R_User(Targ8.RUSER),
        .Targ8_Aw_Lock(Targ8.AWLOCK),
        .Targ8_Ar_Lock(Targ8.ARLOCK),
        .Targ8_Aw_Id(Targ8.AWID),
        .Targ8_Ar_Len(Targ8.ARLEN),
        .Targ8_Ar_User(Targ8.ARUSER),
        .Targ8_B_Id(Targ8.BID),
        .Targ8_W_Valid(Targ8.WVALID),
        .Targ8_B_Ready(Targ8.BREADY),
        .Targ8_W_Data(Targ8.WDATA),
        .Targ8_R_Valid(Targ8.RVALID),
        .Targ8_R_Data(Targ8.RDATA),
        .Targ8_R_Id(Targ8.RID),
        .Targ8_B_Resp(Targ8.BRESP),
        .Targ8_Aw_Size(Targ8.AWSIZE),
        .Targ8_Aw_Addr(Targ8.AWADDR),
        .Targ8_Aw_Cache(Targ8.AWCACHE),
        .Targ8_W_Last(Targ8.WLAST),
        .Targ8_R_Ready(Targ8.RREADY),
        .Targ8_Ar_Ready(Targ8.ARREADY),
        .Targ8_Ar_Cache(Targ8.ARCACHE),
        .Targ8_R_Last(Targ8.RLAST),
        .Targ8_Aw_Qos(Targ8.AWQOS),
        .Targ8_Ar_Valid(Targ8.ARVALID),
        .Targ8_Aw_User(Targ8.AWUSER),
        .Targ8_Ar_Size(Targ8.ARSIZE),
        .Targ8_Aw_Ready(Targ8.AWREADY),
        .Targ8_W_Id(Targ8.WID),
        .Targ8_B_User(Targ8.BUSER),
        .Targ8_Ar_Prot(Targ8.ARPROT),
        .Targ8_Ar_Burst(Targ8.ARBURST),
        .Targ8_R_Resp(Targ8.RRESP),
        .Targ8_Aw_Len(Targ8.AWLEN),
        .Targ8_Aw_Prot(Targ8.AWPROT),
        .Targ8_W_Strb(Targ8.WSTRB),
        .Targ8_Aw_Burst(Targ8.AWBURST),
        .Targ8_B_Valid(Targ8.BVALID),
        .Targ5_Ar_Addr(Targ5.ARADDR),
        .Targ5_W_Ready(Targ5.WREADY),
        .Targ5_Aw_Valid(Targ5.AWVALID),
        .Targ5_Ar_Qos(Targ5.ARQOS),
        .Targ5_Ar_Id(Targ5.ARID),
        .Targ5_R_User(Targ5.RUSER),
        .Targ5_Aw_Lock(Targ5.AWLOCK),
        .Targ5_Ar_Lock(Targ5.ARLOCK),
        .Targ5_Aw_Id(Targ5.AWID),
        .Targ5_Ar_Len(Targ5.ARLEN),
        .Targ5_Ar_User(Targ5.ARUSER),
        .Targ5_B_Id(Targ5.BID),
        .Targ5_W_Valid(Targ5.WVALID),
        .Targ5_B_Ready(Targ5.BREADY),
        .Targ5_W_Data(Targ5.WDATA),
        .Targ5_R_Valid(Targ5.RVALID),
        .Targ5_R_Data(Targ5.RDATA),
        .Targ5_R_Id(Targ5.RID),
        .Targ5_B_Resp(Targ5.BRESP),
        .Targ5_Aw_Size(Targ5.AWSIZE),
        .Targ5_Aw_Addr(Targ5.AWADDR),
        .Targ5_Aw_Cache(Targ5.AWCACHE),
        .Targ5_W_Last(Targ5.WLAST),
        .Targ5_R_Ready(Targ5.RREADY),
        .Targ5_Ar_Ready(Targ5.ARREADY),
        .Targ5_Ar_Cache(Targ5.ARCACHE),
        .Targ5_R_Last(Targ5.RLAST),
        .Targ5_Aw_Qos(Targ5.AWQOS),
        .Targ5_Ar_Valid(Targ5.ARVALID),
        .Targ5_Aw_User(Targ5.AWUSER),
        .Targ5_Ar_Size(Targ5.ARSIZE),
        .Targ5_Aw_Ready(Targ5.AWREADY),
        .Targ5_W_Id(Targ5.WID),
        .Targ5_B_User(Targ5.BUSER),
        .Targ5_Ar_Prot(Targ5.ARPROT),
        .Targ5_Ar_Burst(Targ5.ARBURST),
        .Targ5_R_Resp(Targ5.RRESP),
        .Targ5_Aw_Len(Targ5.AWLEN),
        .Targ5_Aw_Prot(Targ5.AWPROT),
        .Targ5_W_Strb(Targ5.WSTRB),
        .Targ5_Aw_Burst(Targ5.AWBURST),
        .Targ5_B_Valid(Targ5.BVALID),
        .Targ4_Ar_Addr(Targ4.ARADDR),
        .Targ4_W_Ready(Targ4.WREADY),
        .Targ4_Aw_Valid(Targ4.AWVALID),
        .Targ4_Ar_Qos(Targ4.ARQOS),
        .Targ4_Ar_Id(Targ4.ARID),
        .Targ4_R_User(Targ4.RUSER),
        .Targ4_Aw_Lock(Targ4.AWLOCK),
        .Targ4_Ar_Lock(Targ4.ARLOCK),
        .Targ4_Aw_Id(Targ4.AWID),
        .Targ4_Ar_Len(Targ4.ARLEN),
        .Targ4_Ar_User(Targ4.ARUSER),
        .Targ4_B_Id(Targ4.BID),
        .Targ4_W_Valid(Targ4.WVALID),
        .Targ4_B_Ready(Targ4.BREADY),
        .Targ4_W_Data(Targ4.WDATA),
        .Targ4_R_Valid(Targ4.RVALID),
        .Targ4_R_Data(Targ4.RDATA),
        .Targ4_R_Id(Targ4.RID),
        .Targ4_B_Resp(Targ4.BRESP),
        .Targ4_Aw_Size(Targ4.AWSIZE),
        .Targ4_Aw_Addr(Targ4.AWADDR),
        .Targ4_Aw_Cache(Targ4.AWCACHE),
        .Targ4_W_Last(Targ4.WLAST),
        .Targ4_R_Ready(Targ4.RREADY),
        .Targ4_Ar_Ready(Targ4.ARREADY),
        .Targ4_Ar_Cache(Targ4.ARCACHE),
        .Targ4_R_Last(Targ4.RLAST),
        .Targ4_Aw_Qos(Targ4.AWQOS),
        .Targ4_Ar_Valid(Targ4.ARVALID),
        .Targ4_Aw_User(Targ4.AWUSER),
        .Targ4_Ar_Size(Targ4.ARSIZE),
        .Targ4_Aw_Ready(Targ4.AWREADY),
        .Targ4_W_Id(Targ4.WID),
        .Targ4_B_User(Targ4.BUSER),
        .Targ4_Ar_Prot(Targ4.ARPROT),
        .Targ4_Ar_Burst(Targ4.ARBURST),
        .Targ4_R_Resp(Targ4.RRESP),
        .Targ4_Aw_Len(Targ4.AWLEN),
        .Targ4_Aw_Prot(Targ4.AWPROT),
        .Targ4_W_Strb(Targ4.WSTRB),
        .Targ4_Aw_Burst(Targ4.AWBURST),
        .Targ4_B_Valid(Targ4.BVALID),
        .Targ7_Ar_Addr(Targ7.ARADDR),
        .Targ7_W_Ready(Targ7.WREADY),
        .Targ7_Aw_Valid(Targ7.AWVALID),
        .Targ7_Ar_Qos(Targ7.ARQOS),
        .Targ7_Ar_Id(Targ7.ARID),
        .Targ7_R_User(Targ7.RUSER),
        .Targ7_Aw_Lock(Targ7.AWLOCK),
        .Targ7_Ar_Lock(Targ7.ARLOCK),
        .Targ7_Aw_Id(Targ7.AWID),
        .Targ7_Ar_Len(Targ7.ARLEN),
        .Targ7_Ar_User(Targ7.ARUSER),
        .Targ7_B_Id(Targ7.BID),
        .Targ7_W_Valid(Targ7.WVALID),
        .Targ7_B_Ready(Targ7.BREADY),
        .Targ7_W_Data(Targ7.WDATA),
        .Targ7_R_Valid(Targ7.RVALID),
        .Targ7_R_Data(Targ7.RDATA),
        .Targ7_R_Id(Targ7.RID),
        .Targ7_B_Resp(Targ7.BRESP),
        .Targ7_Aw_Size(Targ7.AWSIZE),
        .Targ7_Aw_Addr(Targ7.AWADDR),
        .Targ7_Aw_Cache(Targ7.AWCACHE),
        .Targ7_W_Last(Targ7.WLAST),
        .Targ7_R_Ready(Targ7.RREADY),
        .Targ7_Ar_Ready(Targ7.ARREADY),
        .Targ7_Ar_Cache(Targ7.ARCACHE),
        .Targ7_R_Last(Targ7.RLAST),
        .Targ7_Aw_Qos(Targ7.AWQOS),
        .Targ7_Ar_Valid(Targ7.ARVALID),
        .Targ7_Aw_User(Targ7.AWUSER),
        .Targ7_Ar_Size(Targ7.ARSIZE),
        .Targ7_Aw_Ready(Targ7.AWREADY),
        .Targ7_W_Id(Targ7.WID),
        .Targ7_B_User(Targ7.BUSER),
        .Targ7_Ar_Prot(Targ7.ARPROT),
        .Targ7_Ar_Burst(Targ7.ARBURST),
        .Targ7_R_Resp(Targ7.RRESP),
        .Targ7_Aw_Len(Targ7.AWLEN),
        .Targ7_Aw_Prot(Targ7.AWPROT),
        .Targ7_W_Strb(Targ7.WSTRB),
        .Targ7_Aw_Burst(Targ7.AWBURST),
        .Targ7_B_Valid(Targ7.BVALID),
        .Targ6_Ar_Addr(Targ6.ARADDR),
        .Targ6_W_Ready(Targ6.WREADY),
        .Targ6_Aw_Valid(Targ6.AWVALID),
        .Targ6_Ar_Qos(Targ6.ARQOS),
        .Targ6_Ar_Id(Targ6.ARID),
        .Targ6_R_User(Targ6.RUSER),
        .Targ6_Aw_Lock(Targ6.AWLOCK),
        .Targ6_Ar_Lock(Targ6.ARLOCK),
        .Targ6_Aw_Id(Targ6.AWID),
        .Targ6_Ar_Len(Targ6.ARLEN),
        .Targ6_Ar_User(Targ6.ARUSER),
        .Targ6_B_Id(Targ6.BID),
        .Targ6_W_Valid(Targ6.WVALID),
        .Targ6_B_Ready(Targ6.BREADY),
        .Targ6_W_Data(Targ6.WDATA),
        .Targ6_R_Valid(Targ6.RVALID),
        .Targ6_R_Data(Targ6.RDATA),
        .Targ6_R_Id(Targ6.RID),
        .Targ6_B_Resp(Targ6.BRESP),
        .Targ6_Aw_Size(Targ6.AWSIZE),
        .Targ6_Aw_Addr(Targ6.AWADDR),
        .Targ6_Aw_Cache(Targ6.AWCACHE),
        .Targ6_W_Last(Targ6.WLAST),
        .Targ6_R_Ready(Targ6.RREADY),
        .Targ6_Ar_Ready(Targ6.ARREADY),
        .Targ6_Ar_Cache(Targ6.ARCACHE),
        .Targ6_R_Last(Targ6.RLAST),
        .Targ6_Aw_Qos(Targ6.AWQOS),
        .Targ6_Ar_Valid(Targ6.ARVALID),
        .Targ6_Aw_User(Targ6.AWUSER),
        .Targ6_Ar_Size(Targ6.ARSIZE),
        .Targ6_Aw_Ready(Targ6.AWREADY),
        .Targ6_W_Id(Targ6.WID),
        .Targ6_B_User(Targ6.BUSER),
        .Targ6_Ar_Prot(Targ6.ARPROT),
        .Targ6_Ar_Burst(Targ6.ARBURST),
        .Targ6_R_Resp(Targ6.RRESP),
        .Targ6_Aw_Len(Targ6.AWLEN),
        .Targ6_Aw_Prot(Targ6.AWPROT),
        .Targ6_W_Strb(Targ6.WSTRB),
        .Targ6_Aw_Burst(Targ6.AWBURST),
        .Targ6_B_Valid(Targ6.BVALID),
        .Targ1_Ar_Addr(Targ1.ARADDR),
        .Targ1_W_Ready(Targ1.WREADY),
        .Targ1_Aw_Valid(Targ1.AWVALID),
        .Targ1_Ar_Qos(Targ1.ARQOS),
        .Targ1_Ar_Id(Targ1.ARID),
        .Targ1_R_User(Targ1.RUSER),
        .Targ1_Aw_Lock(Targ1.AWLOCK),
        .Targ1_Ar_Lock(Targ1.ARLOCK),
        .Targ1_Aw_Id(Targ1.AWID),
        .Targ1_Ar_Len(Targ1.ARLEN),
        .Targ1_Ar_User(Targ1.ARUSER),
        .Targ1_B_Id(Targ1.BID),
        .Targ1_W_Valid(Targ1.WVALID),
        .Targ1_B_Ready(Targ1.BREADY),
        .Targ1_W_Data(Targ1.WDATA),
        .Targ1_R_Valid(Targ1.RVALID),
        .Targ1_R_Data(Targ1.RDATA),
        .Targ1_R_Id(Targ1.RID),
        .Targ1_B_Resp(Targ1.BRESP),
        .Targ1_Aw_Size(Targ1.AWSIZE),
        .Targ1_Aw_Addr(Targ1.AWADDR),
        .Targ1_Aw_Cache(Targ1.AWCACHE),
        .Targ1_W_Last(Targ1.WLAST),
        .Targ1_R_Ready(Targ1.RREADY),
        .Targ1_Ar_Ready(Targ1.ARREADY),
        .Targ1_Ar_Cache(Targ1.ARCACHE),
        .Targ1_R_Last(Targ1.RLAST),
        .Targ1_Aw_Qos(Targ1.AWQOS),
        .Targ1_Ar_Valid(Targ1.ARVALID),
        .Targ1_Aw_User(Targ1.AWUSER),
        .Targ1_Ar_Size(Targ1.ARSIZE),
        .Targ1_Aw_Ready(Targ1.AWREADY),
        .Targ1_W_Id(Targ1.WID),
        .Targ1_B_User(Targ1.BUSER),
        .Targ1_Ar_Prot(Targ1.ARPROT),
        .Targ1_Ar_Burst(Targ1.ARBURST),
        .Targ1_R_Resp(Targ1.RRESP),
        .Targ1_Aw_Len(Targ1.AWLEN),
        .Targ1_Aw_Prot(Targ1.AWPROT),
        .Targ1_W_Strb(Targ1.WSTRB),
        .Targ1_Aw_Burst(Targ1.AWBURST),
        .Targ1_B_Valid(Targ1.BVALID),
        .Targ0_Ar_Addr(Targ0.ARADDR),
        .Targ0_W_Ready(Targ0.WREADY),
        .Targ0_Aw_Valid(Targ0.AWVALID),
        .Targ0_Ar_Qos(Targ0.ARQOS),
        .Targ0_Ar_Id(Targ0.ARID),
        .Targ0_R_User(Targ0.RUSER),
        .Targ0_Aw_Lock(Targ0.AWLOCK),
        .Targ0_Ar_Lock(Targ0.ARLOCK),
        .Targ0_Aw_Id(Targ0.AWID),
        .Targ0_Ar_Len(Targ0.ARLEN),
        .Targ0_Ar_User(Targ0.ARUSER),
        .Targ0_B_Id(Targ0.BID),
        .Targ0_W_Valid(Targ0.WVALID),
        .Targ0_B_Ready(Targ0.BREADY),
        .Targ0_W_Data(Targ0.WDATA),
        .Targ0_R_Valid(Targ0.RVALID),
        .Targ0_R_Data(Targ0.RDATA),
        .Targ0_R_Id(Targ0.RID),
        .Targ0_B_Resp(Targ0.BRESP),
        .Targ0_Aw_Size(Targ0.AWSIZE),
        .Targ0_Aw_Addr(Targ0.AWADDR),
        .Targ0_Aw_Cache(Targ0.AWCACHE),
        .Targ0_W_Last(Targ0.WLAST),
        .Targ0_R_Ready(Targ0.RREADY),
        .Targ0_Ar_Ready(Targ0.ARREADY),
        .Targ0_Ar_Cache(Targ0.ARCACHE),
        .Targ0_R_Last(Targ0.RLAST),
        .Targ0_Aw_Qos(Targ0.AWQOS),
        .Targ0_Ar_Valid(Targ0.ARVALID),
        .Targ0_Aw_User(Targ0.AWUSER),
        .Targ0_Ar_Size(Targ0.ARSIZE),
        .Targ0_Aw_Ready(Targ0.AWREADY),
        .Targ0_W_Id(Targ0.WID),
        .Targ0_B_User(Targ0.BUSER),
        .Targ0_Ar_Prot(Targ0.ARPROT),
        .Targ0_Ar_Burst(Targ0.ARBURST),
        .Targ0_R_Resp(Targ0.RRESP),
        .Targ0_Aw_Len(Targ0.AWLEN),
        .Targ0_Aw_Prot(Targ0.AWPROT),
        .Targ0_W_Strb(Targ0.WSTRB),
        .Targ0_Aw_Burst(Targ0.AWBURST),
        .Targ0_B_Valid(Targ0.BVALID),
        .Targ3_Ar_Addr(Targ3.ARADDR),
        .Targ3_W_Ready(Targ3.WREADY),
        .Targ3_Aw_Valid(Targ3.AWVALID),
        .Targ3_Ar_Qos(Targ3.ARQOS),
        .Targ3_Ar_Id(Targ3.ARID),
        .Targ3_R_User(Targ3.RUSER),
        .Targ3_Aw_Lock(Targ3.AWLOCK),
        .Targ3_Ar_Lock(Targ3.ARLOCK),
        .Targ3_Aw_Id(Targ3.AWID),
        .Targ3_Ar_Len(Targ3.ARLEN),
        .Targ3_Ar_User(Targ3.ARUSER),
        .Targ3_B_Id(Targ3.BID),
        .Targ3_W_Valid(Targ3.WVALID),
        .Targ3_B_Ready(Targ3.BREADY),
        .Targ3_W_Data(Targ3.WDATA),
        .Targ3_R_Valid(Targ3.RVALID),
        .Targ3_R_Data(Targ3.RDATA),
        .Targ3_R_Id(Targ3.RID),
        .Targ3_B_Resp(Targ3.BRESP),
        .Targ3_Aw_Size(Targ3.AWSIZE),
        .Targ3_Aw_Addr(Targ3.AWADDR),
        .Targ3_Aw_Cache(Targ3.AWCACHE),
        .Targ3_W_Last(Targ3.WLAST),
        .Targ3_R_Ready(Targ3.RREADY),
        .Targ3_Ar_Ready(Targ3.ARREADY),
        .Targ3_Ar_Cache(Targ3.ARCACHE),
        .Targ3_R_Last(Targ3.RLAST),
        .Targ3_Aw_Qos(Targ3.AWQOS),
        .Targ3_Ar_Valid(Targ3.ARVALID),
        .Targ3_Aw_User(Targ3.AWUSER),
        .Targ3_Ar_Size(Targ3.ARSIZE),
        .Targ3_Aw_Ready(Targ3.AWREADY),
        .Targ3_W_Id(Targ3.WID),
        .Targ3_B_User(Targ3.BUSER),
        .Targ3_Ar_Prot(Targ3.ARPROT),
        .Targ3_Ar_Burst(Targ3.ARBURST),
        .Targ3_R_Resp(Targ3.RRESP),
        .Targ3_Aw_Len(Targ3.AWLEN),
        .Targ3_Aw_Prot(Targ3.AWPROT),
        .Targ3_W_Strb(Targ3.WSTRB),
        .Targ3_Aw_Burst(Targ3.AWBURST),
        .Targ3_B_Valid(Targ3.BVALID),
        .Targ2_Ar_Addr(Targ2.ARADDR),
        .Targ2_W_Ready(Targ2.WREADY),
        .Targ2_Aw_Valid(Targ2.AWVALID),
        .Targ2_Ar_Qos(Targ2.ARQOS),
        .Targ2_Ar_Id(Targ2.ARID),
        .Targ2_R_User(Targ2.RUSER),
        .Targ2_Aw_Lock(Targ2.AWLOCK),
        .Targ2_Ar_Lock(Targ2.ARLOCK),
        .Targ2_Aw_Id(Targ2.AWID),
        .Targ2_Ar_Len(Targ2.ARLEN),
        .Targ2_Ar_User(Targ2.ARUSER),
        .Targ2_B_Id(Targ2.BID),
        .Targ2_W_Valid(Targ2.WVALID),
        .Targ2_B_Ready(Targ2.BREADY),
        .Targ2_W_Data(Targ2.WDATA),
        .Targ2_R_Valid(Targ2.RVALID),
        .Targ2_R_Data(Targ2.RDATA),
        .Targ2_R_Id(Targ2.RID),
        .Targ2_B_Resp(Targ2.BRESP),
        .Targ2_Aw_Size(Targ2.AWSIZE),
        .Targ2_Aw_Addr(Targ2.AWADDR),
        .Targ2_Aw_Cache(Targ2.AWCACHE),
        .Targ2_W_Last(Targ2.WLAST),
        .Targ2_R_Ready(Targ2.RREADY),
        .Targ2_Ar_Ready(Targ2.ARREADY),
        .Targ2_Ar_Cache(Targ2.ARCACHE),
        .Targ2_R_Last(Targ2.RLAST),
        .Targ2_Aw_Qos(Targ2.AWQOS),
        .Targ2_Ar_Valid(Targ2.ARVALID),
        .Targ2_Aw_User(Targ2.AWUSER),
        .Targ2_Ar_Size(Targ2.ARSIZE),
        .Targ2_Aw_Ready(Targ2.AWREADY),
        .Targ2_W_Id(Targ2.WID),
        .Targ2_B_User(Targ2.BUSER),
        .Targ2_Ar_Prot(Targ2.ARPROT),
        .Targ2_Ar_Burst(Targ2.ARBURST),
        .Targ2_R_Resp(Targ2.RRESP),
        .Targ2_Aw_Len(Targ2.AWLEN),
        .Targ2_Aw_Prot(Targ2.AWPROT),
        .Targ2_W_Strb(Targ2.WSTRB),
        .Targ2_Aw_Burst(Targ2.AWBURST),
        .Targ2_B_Valid(Targ2.BVALID),
        .Targ11_Ar_Addr(Targ11.ARADDR),
        .Targ11_W_Ready(Targ11.WREADY),
        .Targ11_Aw_Valid(Targ11.AWVALID),
        .Targ11_Ar_Qos(Targ11.ARQOS),
        .Targ11_Ar_Id(Targ11.ARID),
        .Targ11_R_User(Targ11.RUSER),
        .Targ11_Aw_Lock(Targ11.AWLOCK),
        .Targ11_Ar_Lock(Targ11.ARLOCK),
        .Targ11_Aw_Id(Targ11.AWID),
        .Targ11_Ar_Len(Targ11.ARLEN),
        .Targ11_Ar_User(Targ11.ARUSER),
        .Targ11_B_Id(Targ11.BID),
        .Targ11_W_Valid(Targ11.WVALID),
        .Targ11_B_Ready(Targ11.BREADY),
        .Targ11_W_Data(Targ11.WDATA),
        .Targ11_R_Valid(Targ11.RVALID),
        .Targ11_R_Data(Targ11.RDATA),
        .Targ11_R_Id(Targ11.RID),
        .Targ11_B_Resp(Targ11.BRESP),
        .Targ11_Aw_Size(Targ11.AWSIZE),
        .Targ11_Aw_Addr(Targ11.AWADDR),
        .Targ11_Aw_Cache(Targ11.AWCACHE),
        .Targ11_W_Last(Targ11.WLAST),
        .Targ11_R_Ready(Targ11.RREADY),
        .Targ11_Ar_Ready(Targ11.ARREADY),
        .Targ11_Ar_Cache(Targ11.ARCACHE),
        .Targ11_R_Last(Targ11.RLAST),
        .Targ11_Aw_Qos(Targ11.AWQOS),
        .Targ11_Ar_Valid(Targ11.ARVALID),
        .Targ11_Aw_User(Targ11.AWUSER),
        .Targ11_Ar_Size(Targ11.ARSIZE),
        .Targ11_Aw_Ready(Targ11.AWREADY),
        .Targ11_W_Id(Targ11.WID),
        .Targ11_B_User(Targ11.BUSER),
        .Targ11_Ar_Prot(Targ11.ARPROT),
        .Targ11_Ar_Burst(Targ11.ARBURST),
        .Targ11_R_Resp(Targ11.RRESP),
        .Targ11_Aw_Len(Targ11.AWLEN),
        .Targ11_Aw_Prot(Targ11.AWPROT),
        .Targ11_W_Strb(Targ11.WSTRB),
        .Targ11_Aw_Burst(Targ11.AWBURST),
        .Targ11_B_Valid(Targ11.BVALID),
        .Targ10_Ar_Addr(Targ10.ARADDR),
        .Targ10_W_Ready(Targ10.WREADY),
        .Targ10_Aw_Valid(Targ10.AWVALID),
        .Targ10_Ar_Qos(Targ10.ARQOS),
        .Targ10_Ar_Id(Targ10.ARID),
        .Targ10_R_User(Targ10.RUSER),
        .Targ10_Aw_Lock(Targ10.AWLOCK),
        .Targ10_Ar_Lock(Targ10.ARLOCK),
        .Targ10_Aw_Id(Targ10.AWID),
        .Targ10_Ar_Len(Targ10.ARLEN),
        .Targ10_Ar_User(Targ10.ARUSER),
        .Targ10_B_Id(Targ10.BID),
        .Targ10_W_Valid(Targ10.WVALID),
        .Targ10_B_Ready(Targ10.BREADY),
        .Targ10_W_Data(Targ10.WDATA),
        .Targ10_R_Valid(Targ10.RVALID),
        .Targ10_R_Data(Targ10.RDATA),
        .Targ10_R_Id(Targ10.RID),
        .Targ10_B_Resp(Targ10.BRESP),
        .Targ10_Aw_Size(Targ10.AWSIZE),
        .Targ10_Aw_Addr(Targ10.AWADDR),
        .Targ10_Aw_Cache(Targ10.AWCACHE),
        .Targ10_W_Last(Targ10.WLAST),
        .Targ10_R_Ready(Targ10.RREADY),
        .Targ10_Ar_Ready(Targ10.ARREADY),
        .Targ10_Ar_Cache(Targ10.ARCACHE),
        .Targ10_R_Last(Targ10.RLAST),
        .Targ10_Aw_Qos(Targ10.AWQOS),
        .Targ10_Ar_Valid(Targ10.ARVALID),
        .Targ10_Aw_User(Targ10.AWUSER),
        .Targ10_Ar_Size(Targ10.ARSIZE),
        .Targ10_Aw_Ready(Targ10.AWREADY),
        .Targ10_W_Id(Targ10.WID),
        .Targ10_B_User(Targ10.BUSER),
        .Targ10_Ar_Prot(Targ10.ARPROT),
        .Targ10_Ar_Burst(Targ10.ARBURST),
        .Targ10_R_Resp(Targ10.RRESP),
        .Targ10_Aw_Len(Targ10.AWLEN),
        .Targ10_Aw_Prot(Targ10.AWPROT),
        .Targ10_W_Strb(Targ10.WSTRB),
        .Targ10_Aw_Burst(Targ10.AWBURST),
        .Targ10_B_Valid(Targ10.BVALID),
        .tm(unbound)        
      );


endmodule
/* verilator lint_on WIDTH */        

