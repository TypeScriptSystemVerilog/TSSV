
        

        
/* verilator lint_off WIDTH */        
module AXI4XBar2x4 
   (
   input logic  clk
   );

   



endmodule
/* verilator lint_on WIDTH */        
